
module signed_mult5760 (out, a, b);

  output     [17:0]  out;
  input   signed  [17:0]   a;
  input   signed  [17:0]   b;
  
  wire  signed  [17:0]  out;
  wire   signed  [35:0]  mult_out;

  assign mult_out = a * b;
  //assign out = mult_out[33:17];
  assign out = {mult_out[35], mult_out[32:16]};
endmodule
