module testVect (
output reg signed [15:0] aud [0:1999]
);

initial begin
aud[0]=16'hf09;
aud[1]=16'h683c;
aud[2]=16'h6199;
aud[3]=16'h13b;
aud[4]=16'h9fbc;
aud[5]=16'h96be;
aud[6]=16'hee86;
aud[7]=16'h5660;
aud[8]=16'h6ed0;
aud[9]=16'h215f;
aud[10]=16'hb540;
aud[11]=16'h8dda;
aud[12]=16'hcf68;
aud[13]=16'h3da2;
aud[14]=16'h7333;
aud[15]=16'h3ed9;
aud[16]=16'hd0b8;
aud[17]=16'h8e0f;
aud[18]=16'hb428;
aud[19]=16'h1ffc;
aud[20]=16'h6e68;
aud[21]=16'h5752;
aud[22]=16'heff4;
aud[23]=16'h9756;
aud[24]=16'h9ef3;
aud[25]=16'hffca;
aud[26]=16'h60d3;
aud[27]=16'h68d7;
aud[28]=16'h1078;
aud[29]=16'ha8f5;
aud[30]=16'h9179;
aud[31]=16'hdf9c;
aud[32]=16'h4b86;
aud[33]=16'h7201;
aud[34]=16'h2fab;
aud[35]=16'hc182;
aud[36]=16'h8ccd;
aud[37]=16'hc202;
aud[38]=16'h3036;
aud[39]=16'h7217;
aud[40]=16'h4b13;
aud[41]=16'hdf09;
aud[42]=16'h914e;
aud[43]=16'ha959;
aud[44]=16'h110e;
aud[45]=16'h6916;
aud[46]=16'h6080;
aud[47]=16'hff31;
aud[48]=16'h9ea1;
aud[49]=16'h9796;
aud[50]=16'hf08b;
aud[51]=16'h57b6;
aud[52]=16'h6e3c;
aud[53]=16'h1f6a;
aud[54]=16'hb3b5;
aud[55]=16'h8e25;
aud[56]=16'hd143;
aud[57]=16'h3f59;
aud[58]=16'h7331;
aud[59]=16'h3d21;
aud[60]=16'hcedd;
aud[61]=16'h8dc6;
aud[62]=16'hb5b4;
aud[63]=16'h21f0;
aud[64]=16'h6ef9;
aud[65]=16'h55fa;
aud[66]=16'hedf0;
aud[67]=16'h9680;
aud[68]=16'ha010;
aud[69]=16'h1d4;
aud[70]=16'h61ea;
aud[71]=16'h67fa;
aud[72]=16'he72;
aud[73]=16'ha7a2;
aud[74]=16'h9210;
aud[75]=16'he192;
aud[76]=16'h4d0e;
aud[77]=16'h71b2;
aud[78]=16'h2dce;
aud[79]=16'hbfce;
aud[80]=16'h8cd3;
aud[81]=16'hc3bd;
aud[82]=16'h320e;
aud[83]=16'h725a;
aud[84]=16'h4984;
aud[85]=16'hdd17;
aud[86]=16'h90c2;
aud[87]=16'haab4;
aud[88]=16'h1312;
aud[89]=16'h69e7;
aud[90]=16'h5f5f;
aud[91]=16'hfd27;
aud[92]=16'h9d8e;
aud[93]=16'h9877;
aud[94]=16'hf291;
aud[95]=16'h5905;
aud[96]=16'h6da0;
aud[97]=16'h1d72;
aud[98]=16'hb231;
aud[99]=16'h8e7a;
aud[100]=16'hd322;
aud[101]=16'h410a;
aud[102]=16'h7327;
aud[103]=16'h3b64;
aud[104]=16'hcd07;
aud[105]=16'h8d87;
aud[106]=16'hb746;
aud[107]=16'h23e2;
aud[108]=16'h6f81;
aud[109]=16'h549c;
aud[110]=16'hebed;
aud[111]=16'h95b3;
aud[112]=16'ha135;
aud[113]=16'h3de;
aud[114]=16'h62f9;
aud[115]=16'h6715;
aud[116]=16'hc6c;
aud[117]=16'ha657;
aud[118]=16'h92b1;
aud[119]=16'he38b;
aud[120]=16'h4e8f;
aud[121]=16'h7159;
aud[122]=16'h2bed;
aud[123]=16'hbe1f;
aud[124]=16'h8ce2;
aud[125]=16'hc57c;
aud[126]=16'h33e2;
aud[127]=16'h7295;
aud[128]=16'h47ef;
aud[129]=16'hdb26;
aud[130]=16'h903f;
aud[131]=16'hac16;
aud[132]=16'h1514;
aud[133]=16'h6ab1;
aud[134]=16'h5e36;
aud[135]=16'hfb1d;
aud[136]=16'h9c83;
aud[137]=16'h9960;
aud[138]=16'hf498;
aud[139]=16'h5a4c;
aud[140]=16'h6cfc;
aud[141]=16'h1b78;
aud[142]=16'hb0b3;
aud[143]=16'h8ed7;
aud[144]=16'hd504;
aud[145]=16'h42b7;
aud[146]=16'h7313;
aud[147]=16'h39a3;
aud[148]=16'hcb35;
aud[149]=16'h8d51;
aud[150]=16'hb8dd;
aud[151]=16'h25d1;
aud[152]=16'h6fff;
aud[153]=16'h5336;
aud[154]=16'he9ec;
aud[155]=16'h94ee;
aud[156]=16'ha261;
aud[157]=16'h5e7;
aud[158]=16'h6400;
aud[159]=16'h6628;
aud[160]=16'ha64;
aud[161]=16'ha512;
aud[162]=16'h935a;
aud[163]=16'he586;
aud[164]=16'h5009;
aud[165]=16'h70f7;
aud[166]=16'h2a09;
aud[167]=16'hbc75;
aud[168]=16'h8cfb;
aud[169]=16'hc740;
aud[170]=16'h35b2;
aud[171]=16'h72c6;
aud[172]=16'h4654;
aud[173]=16'hd939;
aud[174]=16'h8fc5;
aud[175]=16'had7f;
aud[176]=16'h1714;
aud[177]=16'h6b71;
aud[178]=16'h5d06;
aud[179]=16'hf914;
aud[180]=16'h9b7f;
aud[181]=16'h9a52;
aud[182]=16'hf6a0;
aud[183]=16'h5b8d;
aud[184]=16'h6c4e;
aud[185]=16'h197c;
aud[186]=16'haf3c;
aud[187]=16'h8f3d;
aud[188]=16'hd6eb;
aud[189]=16'h445e;
aud[190]=16'h72f6;
aud[191]=16'h37dc;
aud[192]=16'hc967;
aud[193]=16'h8d24;
aud[194]=16'hba7b;
aud[195]=16'h27bc;
aud[196]=16'h7075;
aud[197]=16'h51c9;
aud[198]=16'he7ec;
aud[199]=16'h9432;
aud[200]=16'ha395;
aud[201]=16'h7f0;
aud[202]=16'h64ff;
aud[203]=16'h6533;
aud[204]=16'h85c;
aud[205]=16'ha3d6;
aud[206]=16'h940c;
aud[207]=16'he783;
aud[208]=16'h517d;
aud[209]=16'h708c;
aud[210]=16'h2821;
aud[211]=16'hbad1;
aud[212]=16'h8d1c;
aud[213]=16'hc908;
aud[214]=16'h377e;
aud[215]=16'h72ef;
aud[216]=16'h44b4;
aud[217]=16'hd74f;
aud[218]=16'h8f53;
aud[219]=16'haeef;
aud[220]=16'h1913;
aud[221]=16'h6c29;
aud[222]=16'h5bce;
aud[223]=16'hf70b;
aud[224]=16'h9a84;
aud[225]=16'h9b4b;
aud[226]=16'hf8a9;
aud[227]=16'h5cc6;
aud[228]=16'h6b98;
aud[229]=16'h177e;
aud[230]=16'hadcb;
aud[231]=16'h8fad;
aud[232]=16'hd8d4;
aud[233]=16'h45ff;
aud[234]=16'h72d0;
aud[235]=16'h3612;
aud[236]=16'hc79e;
aud[237]=16'h8d01;
aud[238]=16'hbc1e;
aud[239]=16'h29a5;
aud[240]=16'h70e2;
aud[241]=16'h5057;
aud[242]=16'he5ee;
aud[243]=16'h937e;
aud[244]=16'ha4d0;
aud[245]=16'h9f9;
aud[246]=16'h65f6;
aud[247]=16'h6435;
aud[248]=16'h653;
aud[249]=16'ha2a0;
aud[250]=16'h94c6;
aud[251]=16'he982;
aud[252]=16'h52eb;
aud[253]=16'h7018;
aud[254]=16'h2636;
aud[255]=16'hb932;
aud[256]=16'h8d47;
aud[257]=16'hcad5;
aud[258]=16'h3945;
aud[259]=16'h730e;
aud[260]=16'h430e;
aud[261]=16'hd568;
aud[262]=16'h8eeb;
aud[263]=16'hb065;
aud[264]=16'h1b10;
aud[265]=16'h6cd9;
aud[266]=16'h5a8f;
aud[267]=16'hf503;
aud[268]=16'h9991;
aud[269]=16'h9c4d;
aud[270]=16'hfab2;
aud[271]=16'h5df8;
aud[272]=16'h6ad9;
aud[273]=16'h157e;
aud[274]=16'hac60;
aud[275]=16'h9025;
aud[276]=16'hdac0;
aud[277]=16'h479b;
aud[278]=16'h72a0;
aud[279]=16'h3442;
aud[280]=16'hc5d9;
aud[281]=16'h8ce6;
aud[282]=16'hbdc7;
aud[283]=16'h2b8a;
aud[284]=16'h7145;
aud[285]=16'h4edd;
aud[286]=16'he3f3;
aud[287]=16'h92d3;
aud[288]=16'ha613;
aud[289]=16'hc01;
aud[290]=16'h66e5;
aud[291]=16'h6330;
aud[292]=16'h449;
aud[293]=16'ha172;
aud[294]=16'h958a;
aud[295]=16'heb83;
aud[296]=16'h5452;
aud[297]=16'h6f9c;
aud[298]=16'h2448;
aud[299]=16'hb799;
aud[300]=16'h8d7b;
aud[301]=16'hcca7;
aud[302]=16'h3b08;
aud[303]=16'h7323;
aud[304]=16'h4163;
aud[305]=16'hd385;
aud[306]=16'h8e8c;
aud[307]=16'hb1e2;
aud[308]=16'h1d0a;
aud[309]=16'h6d7f;
aud[310]=16'h5949;
aud[311]=16'hf2fc;
aud[312]=16'h98a7;
aud[313]=16'h9d56;
aud[314]=16'hfcbc;
aud[315]=16'h5f22;
aud[316]=16'h6a12;
aud[317]=16'h137c;
aud[318]=16'haafd;
aud[319]=16'h90a6;
aud[320]=16'hdcb0;
aud[321]=16'h4931;
aud[322]=16'h7267;
aud[323]=16'h326f;
aud[324]=16'hc418;
aud[325]=16'h8cd5;
aud[326]=16'hbf74;
aud[327]=16'h2d6b;
aud[328]=16'h71a0;
aud[329]=16'h4d5d;
aud[330]=16'he1fa;
aud[331]=16'h9231;
aud[332]=16'ha75d;
aud[333]=16'he07;
aud[334]=16'h67cc;
aud[335]=16'h6222;
aud[336]=16'h23f;
aud[337]=16'ha04c;
aud[338]=16'h9655;
aud[339]=16'hed85;
aud[340]=16'h55b3;
aud[341]=16'h6f16;
aud[342]=16'h2257;
aud[343]=16'hb606;
aud[344]=16'h8db8;
aud[345]=16'hce7c;
aud[346]=16'h3cc6;
aud[347]=16'h7330;
aud[348]=16'h3fb3;
aud[349]=16'hd1a5;
aud[350]=16'h8e36;
aud[351]=16'hb365;
aud[352]=16'h1f02;
aud[353]=16'h6e1d;
aud[354]=16'h57fb;
aud[355]=16'hf0f6;
aud[356]=16'h97c4;
aud[357]=16'h9e68;
aud[358]=16'hfec6;
aud[359]=16'h6045;
aud[360]=16'h6942;
aud[361]=16'h1179;
aud[362]=16'ha9a0;
aud[363]=16'h9131;
aud[364]=16'hdea2;
aud[365]=16'h4ac1;
aud[366]=16'h7225;
aud[367]=16'h3098;
aud[368]=16'hc25d;
aud[369]=16'h8ccd;
aud[370]=16'hc127;
aud[371]=16'h2f49;
aud[372]=16'h71f2;
aud[373]=16'h4bd8;
aud[374]=16'he003;
aud[375]=16'h9197;
aud[376]=16'ha8ae;
aud[377]=16'h100d;
aud[378]=16'h68aa;
aud[379]=16'h610d;
aud[380]=16'h35;
aud[381]=16'h9f2d;
aud[382]=16'h972a;
aud[383]=16'hef89;
aud[384]=16'h570c;
aud[385]=16'h6e87;
aud[386]=16'h2064;
aud[387]=16'hb479;
aud[388]=16'h8dff;
aud[389]=16'hd055;
aud[390]=16'h3e7f;
aud[391]=16'h7333;
aud[392]=16'h3dfd;
aud[393]=16'hcfc9;
aud[394]=16'h8de9;
aud[395]=16'hb4ee;
aud[396]=16'h20f7;
aud[397]=16'h6eb2;
aud[398]=16'h56a7;
aud[399]=16'heef1;
aud[400]=16'h96ea;
aud[401]=16'h9f81;
aud[402]=16'hd0;
aud[403]=16'h6160;
aud[404]=16'h6869;
aud[405]=16'hf74;
aud[406]=16'ha84a;
aud[407]=16'h91c4;
aud[408]=16'he097;
aud[409]=16'h4c4b;
aud[410]=16'h71da;
aud[411]=16'h2ebc;
aud[412]=16'hc0a6;
aud[413]=16'h8ccf;
aud[414]=16'hc2df;
aud[415]=16'h3123;
aud[416]=16'h723a;
aud[417]=16'h4a4c;
aud[418]=16'hde0f;
aud[419]=16'h9107;
aud[420]=16'haa06;
aud[421]=16'h1211;
aud[422]=16'h6980;
aud[423]=16'h5ff0;
aud[424]=16'hfe2b;
aud[425]=16'h9e16;
aud[426]=16'h9806;
aud[427]=16'hf18f;
aud[428]=16'h585f;
aud[429]=16'h6def;
aud[430]=16'h1e6d;
aud[431]=16'hb2f2;
aud[432]=16'h8e4f;
aud[433]=16'hd233;
aud[434]=16'h4033;
aud[435]=16'h732d;
aud[436]=16'h3c43;
aud[437]=16'hcdf1;
aud[438]=16'h8da5;
aud[439]=16'hb67d;
aud[440]=16'h22ea;
aud[441]=16'h6f3e;
aud[442]=16'h554b;
aud[443]=16'heced;
aud[444]=16'h9618;
aud[445]=16'ha0a2;
aud[446]=16'h2da;
aud[447]=16'h6273;
aud[448]=16'h6788;
aud[449]=16'hd6e;
aud[450]=16'ha6fb;
aud[451]=16'h9260;
aud[452]=16'he28f;
aud[453]=16'h4dcf;
aud[454]=16'h7186;
aud[455]=16'h2cdd;
aud[456]=16'hbef5;
aud[457]=16'h8cd9;
aud[458]=16'hc49c;
aud[459]=16'h32fa;
aud[460]=16'h7279;
aud[461]=16'h48ba;
aud[462]=16'hdc1d;
aud[463]=16'h907f;
aud[464]=16'hab65;
aud[465]=16'h1414;
aud[466]=16'h6a4d;
aud[467]=16'h5ecb;
aud[468]=16'hfc21;
aud[469]=16'h9d07;
aud[470]=16'h98eb;
aud[471]=16'hf395;
aud[472]=16'h59aa;
aud[473]=16'h6d4f;
aud[474]=16'h1c75;
aud[475]=16'hb171;
aud[476]=16'h8ea7;
aud[477]=16'hd414;
aud[478]=16'h41e2;
aud[479]=16'h731e;
aud[480]=16'h3a83;
aud[481]=16'hcc1d;
aud[482]=16'h8d6b;
aud[483]=16'hb812;
aud[484]=16'h24da;
aud[485]=16'h6fc1;
aud[486]=16'h53e9;
aud[487]=16'heaeb;
aud[488]=16'h954f;
aud[489]=16'ha1ca;
aud[490]=16'h4e3;
aud[491]=16'h637e;
aud[492]=16'h669f;
aud[493]=16'hb67;
aud[494]=16'ha5b3;
aud[495]=16'h9305;
aud[496]=16'he489;
aud[497]=16'h4f4d;
aud[498]=16'h7129;
aud[499]=16'h2afb;
aud[500]=16'hbd49;
aud[501]=16'h8ced;
aud[502]=16'hc65e;
aud[503]=16'h34cc;
aud[504]=16'h72af;
aud[505]=16'h4722;
aud[506]=16'hda2f;
aud[507]=16'h9000;
aud[508]=16'haccb;
aud[509]=16'h1615;
aud[510]=16'h6b12;
aud[511]=16'h5d9e;
aud[512]=16'hfa18;
aud[513]=16'h9c00;
aud[514]=16'h99d8;
aud[515]=16'hf59d;
aud[516]=16'h5aee;
aud[517]=16'h6ca6;
aud[518]=16'h1a7a;
aud[519]=16'haff6;
aud[520]=16'h8f09;
aud[521]=16'hd5f8;
aud[522]=16'h438c;
aud[523]=16'h7305;
aud[524]=16'h38bf;
aud[525]=16'hca4d;
aud[526]=16'h8d39;
aud[527]=16'hb9ac;
aud[528]=16'h26c8;
aud[529]=16'h703c;
aud[530]=16'h5280;
aud[531]=16'he8eb;
aud[532]=16'h948e;
aud[533]=16'ha2fb;
aud[534]=16'h6ed;
aud[535]=16'h6481;
aud[536]=16'h65ae;
aud[537]=16'h95f;
aud[538]=16'ha473;
aud[539]=16'h93b2;
aud[540]=16'he685;
aud[541]=16'h50c5;
aud[542]=16'h70c3;
aud[543]=16'h2915;
aud[544]=16'hbba2;
aud[545]=16'h8d0a;
aud[546]=16'hc824;
aud[547]=16'h369a;
aud[548]=16'h72dc;
aud[549]=16'h4584;
aud[550]=16'hd843;
aud[551]=16'h8f8b;
aud[552]=16'hae37;
aud[553]=16'h1815;
aud[554]=16'h6bcf;
aud[555]=16'h5c6a;
aud[556]=16'hf80f;
aud[557]=16'h9b00;
aud[558]=16'h9ace;
aud[559]=16'hf7a5;
aud[560]=16'h5c2b;
aud[561]=16'h6bf4;
aud[562]=16'h187c;
aud[563]=16'hae82;
aud[564]=16'h8f74;
aud[565]=16'hd7e0;
aud[566]=16'h4530;
aud[567]=16'h72e4;
aud[568]=16'h36f7;
aud[569]=16'hc881;
aud[570]=16'h8d11;
aud[571]=16'hbb4d;
aud[572]=16'h28b2;
aud[573]=16'h70ad;
aud[574]=16'h5110;
aud[575]=16'he6ec;
aud[576]=16'h93d6;
aud[577]=16'ha432;
aud[578]=16'h8f6;
aud[579]=16'h657c;
aud[580]=16'h64b5;
aud[581]=16'h757;
aud[582]=16'ha339;
aud[583]=16'h9468;
aud[584]=16'he883;
aud[585]=16'h5236;
aud[586]=16'h7053;
aud[587]=16'h272b;
aud[588]=16'hba00;
aud[589]=16'h8d31;
aud[590]=16'hc9ef;
aud[591]=16'h3863;
aud[592]=16'h72ff;
aud[593]=16'h43e1;
aud[594]=16'hd65b;
aud[595]=16'h8f1e;
aud[596]=16'hafaa;
aud[597]=16'h1a12;
aud[598]=16'h6c82;
aud[599]=16'h5b2f;
aud[600]=16'hf606;
aud[601]=16'h9a09;
aud[602]=16'h9bcb;
aud[603]=16'hf9ae;
aud[604]=16'h5d60;
aud[605]=16'h6b39;
aud[606]=16'h167d;
aud[607]=16'had14;
aud[608]=16'h8fe8;
aud[609]=16'hd9cb;
aud[610]=16'h46ce;
aud[611]=16'h72b9;
aud[612]=16'h352a;
aud[613]=16'hc6ba;
aud[614]=16'h8cf2;
aud[615]=16'hbcf2;
aud[616]=16'h2a98;
aud[617]=16'h7115;
aud[618]=16'h4f9a;
aud[619]=16'he4f0;
aud[620]=16'h9327;
aud[621]=16'ha571;
aud[622]=16'hafe;
aud[623]=16'h666f;
aud[624]=16'h63b3;
aud[625]=16'h54d;
aud[626]=16'ha208;
aud[627]=16'h9527;
aud[628]=16'hea83;
aud[629]=16'h53a0;
aud[630]=16'h6fdb;
aud[631]=16'h253f;
aud[632]=16'hb864;
aud[633]=16'h8d60;
aud[634]=16'hcbbe;
aud[635]=16'h3a28;
aud[636]=16'h731a;
aud[637]=16'h4239;
aud[638]=16'hd476;
aud[639]=16'h8eba;
aud[640]=16'hb123;
aud[641]=16'h1c0e;
aud[642]=16'h6d2d;
aud[643]=16'h59ec;
aud[644]=16'hf3ff;
aud[645]=16'h991b;
aud[646]=16'h9cd1;
aud[647]=16'hfbb8;
aud[648]=16'h5e8e;
aud[649]=16'h6a76;
aud[650]=16'h147c;
aud[651]=16'habad;
aud[652]=16'h9065;
aud[653]=16'hdbb9;
aud[654]=16'h4867;
aud[655]=16'h7285;
aud[656]=16'h3358;
aud[657]=16'hc4f7;
aud[658]=16'h8cdd;
aud[659]=16'hbe9e;
aud[660]=16'h2c7c;
aud[661]=16'h7174;
aud[662]=16'h4e1d;
aud[663]=16'he2f5;
aud[664]=16'h9281;
aud[665]=16'ha6b8;
aud[666]=16'hd05;
aud[667]=16'h675a;
aud[668]=16'h62a9;
aud[669]=16'h344;
aud[670]=16'ha0dd;
aud[671]=16'h95ef;
aud[672]=16'hec85;
aud[673]=16'h5504;
aud[674]=16'h6f59;
aud[675]=16'h234f;
aud[676]=16'hb6ce;
aud[677]=16'h8d99;
aud[678]=16'hcd92;
aud[679]=16'h3be8;
aud[680]=16'h732b;
aud[681]=16'h408b;
aud[682]=16'hd294;
aud[683]=16'h8e60;
aud[684]=16'hb2a3;
aud[685]=16'h1e07;
aud[686]=16'h6dcf;
aud[687]=16'h58a2;
aud[688]=16'hf1f8;
aud[689]=16'h9834;
aud[690]=16'h9dde;
aud[691]=16'hfdc1;
aud[692]=16'h5fb5;
aud[693]=16'h69aa;
aud[694]=16'h127a;
aud[695]=16'haa4d;
aud[696]=16'h90eb;
aud[697]=16'hddaa;
aud[698]=16'h49fa;
aud[699]=16'h7247;
aud[700]=16'h3183;
aud[701]=16'hc339;
aud[702]=16'h8cd0;
aud[703]=16'hc04e;
aud[704]=16'h2e5b;
aud[705]=16'h71ca;
aud[706]=16'h4c9b;
aud[707]=16'he0fd;
aud[708]=16'h91e3;
aud[709]=16'ha805;
aud[710]=16'hf0b;
aud[711]=16'h683c;
aud[712]=16'h6198;
aud[713]=16'h13a;
aud[714]=16'h9fbb;
aud[715]=16'h96bf;
aud[716]=16'hee88;
aud[717]=16'h5661;
aud[718]=16'h6ecf;
aud[719]=16'h215d;
aud[720]=16'hb53e;
aud[721]=16'h8ddb;
aud[722]=16'hcf69;
aud[723]=16'h3da4;
aud[724]=16'h7333;
aud[725]=16'h3ed8;
aud[726]=16'hd0b6;
aud[727]=16'h8e0e;
aud[728]=16'hb429;
aud[729]=16'h1ffe;
aud[730]=16'h6e69;
aud[731]=16'h5751;
aud[732]=16'heff2;
aud[733]=16'h9756;
aud[734]=16'h9ef4;
aud[735]=16'hffcb;
aud[736]=16'h60d4;
aud[737]=16'h68d6;
aud[738]=16'h1076;
aud[739]=16'ha8f3;
aud[740]=16'h9179;
aud[741]=16'hdf9d;
aud[742]=16'h4b88;
aud[743]=16'h7201;
aud[744]=16'h2faa;
aud[745]=16'hc180;
aud[746]=16'h8ccd;
aud[747]=16'hc204;
aud[748]=16'h3038;
aud[749]=16'h7217;
aud[750]=16'h4b12;
aud[751]=16'hdf08;
aud[752]=16'h914e;
aud[753]=16'ha95a;
aud[754]=16'h1110;
aud[755]=16'h6916;
aud[756]=16'h607f;
aud[757]=16'hff2f;
aud[758]=16'h9ea0;
aud[759]=16'h9797;
aud[760]=16'hf08d;
aud[761]=16'h57b7;
aud[762]=16'h6e3c;
aud[763]=16'h1f68;
aud[764]=16'hb3b4;
aud[765]=16'h8e26;
aud[766]=16'hd144;
aud[767]=16'h3f5a;
aud[768]=16'h7331;
aud[769]=16'h3d20;
aud[770]=16'hcedc;
aud[771]=16'h8dc6;
aud[772]=16'hb5b5;
aud[773]=16'h21f2;
aud[774]=16'h6ef9;
aud[775]=16'h55f9;
aud[776]=16'hedee;
aud[777]=16'h9680;
aud[778]=16'ha011;
aud[779]=16'h1d6;
aud[780]=16'h61eb;
aud[781]=16'h67f9;
aud[782]=16'he70;
aud[783]=16'ha7a1;
aud[784]=16'h9211;
aud[785]=16'he194;
aud[786]=16'h4d0f;
aud[787]=16'h71b1;
aud[788]=16'h2dcd;
aud[789]=16'hbfcc;
aud[790]=16'h8cd3;
aud[791]=16'hc3be;
aud[792]=16'h3210;
aud[793]=16'h725b;
aud[794]=16'h4983;
aud[795]=16'hdd15;
aud[796]=16'h90c2;
aud[797]=16'haab5;
aud[798]=16'h1314;
aud[799]=16'h69e8;
aud[800]=16'h5f5e;
aud[801]=16'hfd25;
aud[802]=16'h9d8d;
aud[803]=16'h9878;
aud[804]=16'hf293;
aud[805]=16'h5906;
aud[806]=16'h6da0;
aud[807]=16'h1d70;
aud[808]=16'hb230;
aud[809]=16'h8e7a;
aud[810]=16'hd323;
aud[811]=16'h410c;
aud[812]=16'h7327;
aud[813]=16'h3b63;
aud[814]=16'hcd06;
aud[815]=16'h8d87;
aud[816]=16'hb747;
aud[817]=16'h23e4;
aud[818]=16'h6f81;
aud[819]=16'h549a;
aud[820]=16'hebeb;
aud[821]=16'h95b2;
aud[822]=16'ha136;
aud[823]=16'h3df;
aud[824]=16'h62fa;
aud[825]=16'h6715;
aud[826]=16'hc6a;
aud[827]=16'ha656;
aud[828]=16'h92b1;
aud[829]=16'he38c;
aud[830]=16'h4e90;
aud[831]=16'h7159;
aud[832]=16'h2bec;
aud[833]=16'hbe1d;
aud[834]=16'h8ce2;
aud[835]=16'hc57d;
aud[836]=16'h33e4;
aud[837]=16'h7295;
aud[838]=16'h47ee;
aud[839]=16'hdb25;
aud[840]=16'h903e;
aud[841]=16'hac18;
aud[842]=16'h1516;
aud[843]=16'h6ab1;
aud[844]=16'h5e35;
aud[845]=16'hfb1c;
aud[846]=16'h9c82;
aud[847]=16'h9961;
aud[848]=16'hf49a;
aud[849]=16'h5a4d;
aud[850]=16'h6cfb;
aud[851]=16'h1b76;
aud[852]=16'hb0b2;
aud[853]=16'h8ed7;
aud[854]=16'hd506;
aud[855]=16'h42b8;
aud[856]=16'h7313;
aud[857]=16'h39a1;
aud[858]=16'hcb34;
aud[859]=16'h8d51;
aud[860]=16'hb8df;
aud[861]=16'h25d2;
aud[862]=16'h7000;
aud[863]=16'h5335;
aud[864]=16'he9ea;
aud[865]=16'h94ed;
aud[866]=16'ha262;
aud[867]=16'h5e9;
aud[868]=16'h6401;
aud[869]=16'h6627;
aud[870]=16'ha62;
aud[871]=16'ha511;
aud[872]=16'h935b;
aud[873]=16'he587;
aud[874]=16'h500a;
aud[875]=16'h70f7;
aud[876]=16'h2a07;
aud[877]=16'hbc74;
aud[878]=16'h8cfb;
aud[879]=16'hc741;
aud[880]=16'h35b4;
aud[881]=16'h72c7;
aud[882]=16'h4653;
aud[883]=16'hd938;
aud[884]=16'h8fc4;
aud[885]=16'had81;
aud[886]=16'h1716;
aud[887]=16'h6b72;
aud[888]=16'h5d05;
aud[889]=16'hf912;
aud[890]=16'h9b7f;
aud[891]=16'h9a52;
aud[892]=16'hf6a2;
aud[893]=16'h5b8e;
aud[894]=16'h6c4e;
aud[895]=16'h197a;
aud[896]=16'haf3b;
aud[897]=16'h8f3e;
aud[898]=16'hd6ec;
aud[899]=16'h445f;
aud[900]=16'h72f6;
aud[901]=16'h37db;
aud[902]=16'hc966;
aud[903]=16'h8d24;
aud[904]=16'hba7c;
aud[905]=16'h27be;
aud[906]=16'h7075;
aud[907]=16'h51c8;
aud[908]=16'he7ea;
aud[909]=16'h9431;
aud[910]=16'ha396;
aud[911]=16'h7f2;
aud[912]=16'h6500;
aud[913]=16'h6532;
aud[914]=16'h85a;
aud[915]=16'ha3d5;
aud[916]=16'h940d;
aud[917]=16'he784;
aud[918]=16'h517f;
aud[919]=16'h708c;
aud[920]=16'h2820;
aud[921]=16'hbad0;
aud[922]=16'h8d1c;
aud[923]=16'hc90a;
aud[924]=16'h3780;
aud[925]=16'h72ef;
aud[926]=16'h44b3;
aud[927]=16'hd74e;
aud[928]=16'h8f53;
aud[929]=16'haef0;
aud[930]=16'h1915;
aud[931]=16'h6c2a;
aud[932]=16'h5bcd;
aud[933]=16'hf70a;
aud[934]=16'h9a84;
aud[935]=16'h9b4c;
aud[936]=16'hf8aa;
aud[937]=16'h5cc7;
aud[938]=16'h6b97;
aud[939]=16'h177c;
aud[940]=16'hadca;
aud[941]=16'h8fad;
aud[942]=16'hd8d6;
aud[943]=16'h4600;
aud[944]=16'h72cf;
aud[945]=16'h3610;
aud[946]=16'hc79c;
aud[947]=16'h8d01;
aud[948]=16'hbc1f;
aud[949]=16'h29a6;
aud[950]=16'h70e2;
aud[951]=16'h5055;
aud[952]=16'he5ed;
aud[953]=16'h937d;
aud[954]=16'ha4d2;
aud[955]=16'h9fb;
aud[956]=16'h65f7;
aud[957]=16'h6434;
aud[958]=16'h651;
aud[959]=16'ha29f;
aud[960]=16'h94c7;
aud[961]=16'he984;
aud[962]=16'h52ec;
aud[963]=16'h7018;
aud[964]=16'h2635;
aud[965]=16'hb931;
aud[966]=16'h8d47;
aud[967]=16'hcad7;
aud[968]=16'h3947;
aud[969]=16'h730e;
aud[970]=16'h430d;
aud[971]=16'hd567;
aud[972]=16'h8eeb;
aud[973]=16'hb067;
aud[974]=16'h1b11;
aud[975]=16'h6cd9;
aud[976]=16'h5a8e;
aud[977]=16'hf501;
aud[978]=16'h9991;
aud[979]=16'h9c4d;
aud[980]=16'hfab4;
aud[981]=16'h5df9;
aud[982]=16'h6ad8;
aud[983]=16'h157c;
aud[984]=16'hac5f;
aud[985]=16'h9025;
aud[986]=16'hdac2;
aud[987]=16'h479c;
aud[988]=16'h72a0;
aud[989]=16'h3441;
aud[990]=16'hc5d7;
aud[991]=16'h8ce6;
aud[992]=16'hbdc8;
aud[993]=16'h2b8b;
aud[994]=16'h7146;
aud[995]=16'h4edc;
aud[996]=16'he3f1;
aud[997]=16'h92d2;
aud[998]=16'ha614;
aud[999]=16'hc02;
aud[1000]=16'h66e6;
aud[1001]=16'h632f;
aud[1002]=16'h448;
aud[1003]=16'ha171;
aud[1004]=16'h958a;
aud[1005]=16'heb84;
aud[1006]=16'h5454;
aud[1007]=16'h6f9b;
aud[1008]=16'h2447;
aud[1009]=16'hb798;
aud[1010]=16'h8d7b;
aud[1011]=16'hcca8;
aud[1012]=16'h3b0a;
aud[1013]=16'h7323;
aud[1014]=16'h4162;
aud[1015]=16'hd383;
aud[1016]=16'h8e8c;
aud[1017]=16'hb1e3;
aud[1018]=16'h1d0c;
aud[1019]=16'h6d80;
aud[1020]=16'h5948;
aud[1021]=16'hf2fa;
aud[1022]=16'h98a6;
aud[1023]=16'h9d57;
aud[1024]=16'hfcbd;
aud[1025]=16'h5f23;
aud[1026]=16'h6a11;
aud[1027]=16'h137a;
aud[1028]=16'haafb;
aud[1029]=16'h90a7;
aud[1030]=16'hdcb2;
aud[1031]=16'h4932;
aud[1032]=16'h7267;
aud[1033]=16'h326d;
aud[1034]=16'hc417;
aud[1035]=16'h8cd5;
aud[1036]=16'hbf76;
aud[1037]=16'h2d6d;
aud[1038]=16'h71a0;
aud[1039]=16'h4d5c;
aud[1040]=16'he1f8;
aud[1041]=16'h9230;
aud[1042]=16'ha75e;
aud[1043]=16'he09;
aud[1044]=16'h67cc;
aud[1045]=16'h6221;
aud[1046]=16'h23e;
aud[1047]=16'ha04b;
aud[1048]=16'h9656;
aud[1049]=16'hed87;
aud[1050]=16'h55b4;
aud[1051]=16'h6f15;
aud[1052]=16'h2256;
aud[1053]=16'hb605;
aud[1054]=16'h8db9;
aud[1055]=16'hce7e;
aud[1056]=16'h3cc7;
aud[1057]=16'h7330;
aud[1058]=16'h3fb1;
aud[1059]=16'hd1a4;
aud[1060]=16'h8e36;
aud[1061]=16'hb366;
aud[1062]=16'h1f04;
aud[1063]=16'h6e1e;
aud[1064]=16'h57fa;
aud[1065]=16'hf0f4;
aud[1066]=16'h97c3;
aud[1067]=16'h9e68;
aud[1068]=16'hfec7;
aud[1069]=16'h6046;
aud[1070]=16'h6941;
aud[1071]=16'h1177;
aud[1072]=16'ha99f;
aud[1073]=16'h9131;
aud[1074]=16'hdea4;
aud[1075]=16'h4ac3;
aud[1076]=16'h7225;
aud[1077]=16'h3096;
aud[1078]=16'hc25b;
aud[1079]=16'h8ccd;
aud[1080]=16'hc129;
aud[1081]=16'h2f4b;
aud[1082]=16'h71f2;
aud[1083]=16'h4bd6;
aud[1084]=16'he001;
aud[1085]=16'h9197;
aud[1086]=16'ha8af;
aud[1087]=16'h100f;
aud[1088]=16'h68ab;
aud[1089]=16'h610c;
aud[1090]=16'h34;
aud[1091]=16'h9f2c;
aud[1092]=16'h972a;
aud[1093]=16'hef8b;
aud[1094]=16'h570d;
aud[1095]=16'h6e86;
aud[1096]=16'h2062;
aud[1097]=16'hb478;
aud[1098]=16'h8dff;
aud[1099]=16'hd057;
aud[1100]=16'h3e80;
aud[1101]=16'h7333;
aud[1102]=16'h3dfc;
aud[1103]=16'hcfc8;
aud[1104]=16'h8de9;
aud[1105]=16'hb4ef;
aud[1106]=16'h20f9;
aud[1107]=16'h6eb3;
aud[1108]=16'h56a6;
aud[1109]=16'heeef;
aud[1110]=16'h96e9;
aud[1111]=16'h9f82;
aud[1112]=16'hd1;
aud[1113]=16'h6161;
aud[1114]=16'h6868;
aud[1115]=16'hf72;
aud[1116]=16'ha849;
aud[1117]=16'h91c4;
aud[1118]=16'he099;
aud[1119]=16'h4c4d;
aud[1120]=16'h71da;
aud[1121]=16'h2ebb;
aud[1122]=16'hc0a5;
aud[1123]=16'h8ccf;
aud[1124]=16'hc2e1;
aud[1125]=16'h3125;
aud[1126]=16'h723a;
aud[1127]=16'h4a4a;
aud[1128]=16'hde0d;
aud[1129]=16'h9106;
aud[1130]=16'haa07;
aud[1131]=16'h1213;
aud[1132]=16'h6981;
aud[1133]=16'h5fef;
aud[1134]=16'hfe2a;
aud[1135]=16'h9e15;
aud[1136]=16'h9807;
aud[1137]=16'hf190;
aud[1138]=16'h5860;
aud[1139]=16'h6def;
aud[1140]=16'h1e6c;
aud[1141]=16'hb2f0;
aud[1142]=16'h8e4f;
aud[1143]=16'hd234;
aud[1144]=16'h4035;
aud[1145]=16'h732d;
aud[1146]=16'h3c41;
aud[1147]=16'hcdef;
aud[1148]=16'h8da5;
aud[1149]=16'hb67e;
aud[1150]=16'h22ec;
aud[1151]=16'h6f3f;
aud[1152]=16'h554a;
aud[1153]=16'heceb;
aud[1154]=16'h9618;
aud[1155]=16'ha0a3;
aud[1156]=16'h2db;
aud[1157]=16'h6274;
aud[1158]=16'h6788;
aud[1159]=16'hd6c;
aud[1160]=16'ha6fa;
aud[1161]=16'h9260;
aud[1162]=16'he291;
aud[1163]=16'h4dd1;
aud[1164]=16'h7186;
aud[1165]=16'h2cdc;
aud[1166]=16'hbef3;
aud[1167]=16'h8cd9;
aud[1168]=16'hc49e;
aud[1169]=16'h32fb;
aud[1170]=16'h7279;
aud[1171]=16'h48b8;
aud[1172]=16'hdc1c;
aud[1173]=16'h907f;
aud[1174]=16'hab66;
aud[1175]=16'h1416;
aud[1176]=16'h6a4e;
aud[1177]=16'h5eca;
aud[1178]=16'hfc20;
aud[1179]=16'h9d06;
aud[1180]=16'h98ec;
aud[1181]=16'hf397;
aud[1182]=16'h59ab;
aud[1183]=16'h6d4e;
aud[1184]=16'h1c73;
aud[1185]=16'hb170;
aud[1186]=16'h8ea8;
aud[1187]=16'hd415;
aud[1188]=16'h41e3;
aud[1189]=16'h731e;
aud[1190]=16'h3a82;
aud[1191]=16'hcc1b;
aud[1192]=16'h8d6b;
aud[1193]=16'hb813;
aud[1194]=16'h24dc;
aud[1195]=16'h6fc2;
aud[1196]=16'h53e8;
aud[1197]=16'heae9;
aud[1198]=16'h954e;
aud[1199]=16'ha1cc;
aud[1200]=16'h4e5;
aud[1201]=16'h637f;
aud[1202]=16'h669f;
aud[1203]=16'hb65;
aud[1204]=16'ha5b2;
aud[1205]=16'h9305;
aud[1206]=16'he48a;
aud[1207]=16'h4f4f;
aud[1208]=16'h7129;
aud[1209]=16'h2af9;
aud[1210]=16'hbd47;
aud[1211]=16'h8ced;
aud[1212]=16'hc660;
aud[1213]=16'h34cd;
aud[1214]=16'h72af;
aud[1215]=16'h4720;
aud[1216]=16'hda2d;
aud[1217]=16'h9000;
aud[1218]=16'haccc;
aud[1219]=16'h1617;
aud[1220]=16'h6b13;
aud[1221]=16'h5d9d;
aud[1222]=16'hfa16;
aud[1223]=16'h9bff;
aud[1224]=16'h99d9;
aud[1225]=16'hf59e;
aud[1226]=16'h5aef;
aud[1227]=16'h6ca5;
aud[1228]=16'h1a78;
aud[1229]=16'haff5;
aud[1230]=16'h8f09;
aud[1231]=16'hd5fa;
aud[1232]=16'h438d;
aud[1233]=16'h7305;
aud[1234]=16'h38be;
aud[1235]=16'hca4b;
aud[1236]=16'h8d39;
aud[1237]=16'hb9ae;
aud[1238]=16'h26c9;
aud[1239]=16'h703c;
aud[1240]=16'h527f;
aud[1241]=16'he8e9;
aud[1242]=16'h948e;
aud[1243]=16'ha2fc;
aud[1244]=16'h6ef;
aud[1245]=16'h6482;
aud[1246]=16'h65ad;
aud[1247]=16'h95d;
aud[1248]=16'ha471;
aud[1249]=16'h93b3;
aud[1250]=16'he687;
aud[1251]=16'h50c6;
aud[1252]=16'h70c2;
aud[1253]=16'h2913;
aud[1254]=16'hbba0;
aud[1255]=16'h8d0a;
aud[1256]=16'hc826;
aud[1257]=16'h369b;
aud[1258]=16'h72dc;
aud[1259]=16'h4583;
aud[1260]=16'hd841;
aud[1261]=16'h8f8a;
aud[1262]=16'hae38;
aud[1263]=16'h1817;
aud[1264]=16'h6bcf;
aud[1265]=16'h5c69;
aud[1266]=16'hf80d;
aud[1267]=16'h9b00;
aud[1268]=16'h9acf;
aud[1269]=16'hf7a7;
aud[1270]=16'h5c2c;
aud[1271]=16'h6bf3;
aud[1272]=16'h187b;
aud[1273]=16'hae81;
aud[1274]=16'h8f74;
aud[1275]=16'hd7e1;
aud[1276]=16'h4531;
aud[1277]=16'h72e4;
aud[1278]=16'h36f5;
aud[1279]=16'hc880;
aud[1280]=16'h8d11;
aud[1281]=16'hbb4e;
aud[1282]=16'h28b3;
aud[1283]=16'h70ad;
aud[1284]=16'h510f;
aud[1285]=16'he6ea;
aud[1286]=16'h93d6;
aud[1287]=16'ha433;
aud[1288]=16'h8f7;
aud[1289]=16'h657d;
aud[1290]=16'h64b4;
aud[1291]=16'h755;
aud[1292]=16'ha338;
aud[1293]=16'h9469;
aud[1294]=16'he885;
aud[1295]=16'h5237;
aud[1296]=16'h7053;
aud[1297]=16'h272a;
aud[1298]=16'hb9ff;
aud[1299]=16'h8d31;
aud[1300]=16'hc9f1;
aud[1301]=16'h3865;
aud[1302]=16'h72ff;
aud[1303]=16'h43e0;
aud[1304]=16'hd659;
aud[1305]=16'h8f1e;
aud[1306]=16'hafab;
aud[1307]=16'h1a14;
aud[1308]=16'h6c83;
aud[1309]=16'h5b2e;
aud[1310]=16'hf604;
aud[1311]=16'h9a09;
aud[1312]=16'h9bcc;
aud[1313]=16'hf9b0;
aud[1314]=16'h5d61;
aud[1315]=16'h6b39;
aud[1316]=16'h167c;
aud[1317]=16'had13;
aud[1318]=16'h8fe8;
aud[1319]=16'hd9cc;
aud[1320]=16'h46d0;
aud[1321]=16'h72b9;
aud[1322]=16'h3528;
aud[1323]=16'hc6b8;
aud[1324]=16'h8cf2;
aud[1325]=16'hbcf4;
aud[1326]=16'h2a9a;
aud[1327]=16'h7115;
aud[1328]=16'h4f99;
aud[1329]=16'he4ee;
aud[1330]=16'h9327;
aud[1331]=16'ha573;
aud[1332]=16'haff;
aud[1333]=16'h6670;
aud[1334]=16'h63b2;
aud[1335]=16'h54b;
aud[1336]=16'ha207;
aud[1337]=16'h9528;
aud[1338]=16'hea85;
aud[1339]=16'h53a1;
aud[1340]=16'h6fda;
aud[1341]=16'h253d;
aud[1342]=16'hb863;
aud[1343]=16'h8d60;
aud[1344]=16'hcbc0;
aud[1345]=16'h3a2a;
aud[1346]=16'h731a;
aud[1347]=16'h4237;
aud[1348]=16'hd474;
aud[1349]=16'h8eba;
aud[1350]=16'hb125;
aud[1351]=16'h1c10;
aud[1352]=16'h6d2e;
aud[1353]=16'h59eb;
aud[1354]=16'hf3fd;
aud[1355]=16'h991a;
aud[1356]=16'h9cd2;
aud[1357]=16'hfbb9;
aud[1358]=16'h5e8f;
aud[1359]=16'h6a75;
aud[1360]=16'h147b;
aud[1361]=16'habac;
aud[1362]=16'h9065;
aud[1363]=16'hdbba;
aud[1364]=16'h4869;
aud[1365]=16'h7285;
aud[1366]=16'h3357;
aud[1367]=16'hc4f6;
aud[1368]=16'h8cdd;
aud[1369]=16'hbe9f;
aud[1370]=16'h2c7d;
aud[1371]=16'h7174;
aud[1372]=16'h4e1c;
aud[1373]=16'he2f4;
aud[1374]=16'h9280;
aud[1375]=16'ha6b9;
aud[1376]=16'hd07;
aud[1377]=16'h675b;
aud[1378]=16'h62a9;
aud[1379]=16'h342;
aud[1380]=16'ha0dc;
aud[1381]=16'h95ef;
aud[1382]=16'hec86;
aud[1383]=16'h5505;
aud[1384]=16'h6f59;
aud[1385]=16'h234e;
aud[1386]=16'hb6cd;
aud[1387]=16'h8d99;
aud[1388]=16'hcd93;
aud[1389]=16'h3bea;
aud[1390]=16'h732b;
aud[1391]=16'h4089;
aud[1392]=16'hd292;
aud[1393]=16'h8e5f;
aud[1394]=16'hb2a4;
aud[1395]=16'h1e09;
aud[1396]=16'h6dd0;
aud[1397]=16'h58a1;
aud[1398]=16'hf1f6;
aud[1399]=16'h9833;
aud[1400]=16'h9ddf;
aud[1401]=16'hfdc3;
aud[1402]=16'h5fb6;
aud[1403]=16'h69aa;
aud[1404]=16'h1278;
aud[1405]=16'haa4c;
aud[1406]=16'h90eb;
aud[1407]=16'hddab;
aud[1408]=16'h49fc;
aud[1409]=16'h7247;
aud[1410]=16'h3181;
aud[1411]=16'hc338;
aud[1412]=16'h8cd0;
aud[1413]=16'hc04f;
aud[1414]=16'h2e5d;
aud[1415]=16'h71ca;
aud[1416]=16'h4c99;
aud[1417]=16'he0fc;
aud[1418]=16'h91e2;
aud[1419]=16'ha806;
aud[1420]=16'hf0d;
aud[1421]=16'h683d;
aud[1422]=16'h6197;
aud[1423]=16'h138;
aud[1424]=16'h9fba;
aud[1425]=16'h96bf;
aud[1426]=16'hee8a;
aud[1427]=16'h5662;
aud[1428]=16'h6ecf;
aud[1429]=16'h215b;
aud[1430]=16'hb53d;
aud[1431]=16'h8ddb;
aud[1432]=16'hcf6b;
aud[1433]=16'h3da5;
aud[1434]=16'h7333;
aud[1435]=16'h3ed6;
aud[1436]=16'hd0b4;
aud[1437]=16'h8e0e;
aud[1438]=16'hb42a;
aud[1439]=16'h2000;
aud[1440]=16'h6e69;
aud[1441]=16'h5750;
aud[1442]=16'heff0;
aud[1443]=16'h9755;
aud[1444]=16'h9ef5;
aud[1445]=16'hffcd;
aud[1446]=16'h60d5;
aud[1447]=16'h68d5;
aud[1448]=16'h1074;
aud[1449]=16'ha8f2;
aud[1450]=16'h917a;
aud[1451]=16'hdf9f;
aud[1452]=16'h4b89;
aud[1453]=16'h7201;
aud[1454]=16'h2fa8;
aud[1455]=16'hc17f;
aud[1456]=16'h8ccd;
aud[1457]=16'hc205;
aud[1458]=16'h3039;
aud[1459]=16'h7217;
aud[1460]=16'h4b10;
aud[1461]=16'hdf06;
aud[1462]=16'h914d;
aud[1463]=16'ha95b;
aud[1464]=16'h1112;
aud[1465]=16'h6917;
aud[1466]=16'h607e;
aud[1467]=16'hff2e;
aud[1468]=16'h9e9f;
aud[1469]=16'h9798;
aud[1470]=16'hf08e;
aud[1471]=16'h57b8;
aud[1472]=16'h6e3b;
aud[1473]=16'h1f66;
aud[1474]=16'hb3b3;
aud[1475]=16'h8e26;
aud[1476]=16'hd146;
aud[1477]=16'h3f5c;
aud[1478]=16'h7331;
aud[1479]=16'h3d1e;
aud[1480]=16'hceda;
aud[1481]=16'h8dc6;
aud[1482]=16'hb5b6;
aud[1483]=16'h21f4;
aud[1484]=16'h6efa;
aud[1485]=16'h55f8;
aud[1486]=16'hedec;
aud[1487]=16'h967f;
aud[1488]=16'ha012;
aud[1489]=16'h1d7;
aud[1490]=16'h61eb;
aud[1491]=16'h67f9;
aud[1492]=16'he6f;
aud[1493]=16'ha7a0;
aud[1494]=16'h9211;
aud[1495]=16'he195;
aud[1496]=16'h4d10;
aud[1497]=16'h71b1;
aud[1498]=16'h2dcb;
aud[1499]=16'hbfcb;
aud[1500]=16'h8cd3;
aud[1501]=16'hc3c0;
aud[1502]=16'h3211;
aud[1503]=16'h725b;
aud[1504]=16'h4981;
aud[1505]=16'hdd13;
aud[1506]=16'h90c1;
aud[1507]=16'haab7;
aud[1508]=16'h1315;
aud[1509]=16'h69e9;
aud[1510]=16'h5f5d;
aud[1511]=16'hfd24;
aud[1512]=16'h9d8c;
aud[1513]=16'h9879;
aud[1514]=16'hf294;
aud[1515]=16'h5907;
aud[1516]=16'h6d9f;
aud[1517]=16'h1d6f;
aud[1518]=16'hb22f;
aud[1519]=16'h8e7a;
aud[1520]=16'hd325;
aud[1521]=16'h410d;
aud[1522]=16'h7327;
aud[1523]=16'h3b61;
aud[1524]=16'hcd04;
aud[1525]=16'h8d87;
aud[1526]=16'hb748;
aud[1527]=16'h23e5;
aud[1528]=16'h6f82;
aud[1529]=16'h5499;
aud[1530]=16'hebe9;
aud[1531]=16'h95b2;
aud[1532]=16'ha137;
aud[1533]=16'h3e1;
aud[1534]=16'h62fb;
aud[1535]=16'h6714;
aud[1536]=16'hc68;
aud[1537]=16'ha654;
aud[1538]=16'h92b2;
aud[1539]=16'he38e;
aud[1540]=16'h4e91;
aud[1541]=16'h7158;
aud[1542]=16'h2bea;
aud[1543]=16'hbe1c;
aud[1544]=16'h8ce2;
aud[1545]=16'hc57f;
aud[1546]=16'h33e5;
aud[1547]=16'h7295;
aud[1548]=16'h47ec;
aud[1549]=16'hdb23;
aud[1550]=16'h903e;
aud[1551]=16'hac19;
aud[1552]=16'h1518;
aud[1553]=16'h6ab2;
aud[1554]=16'h5e34;
aud[1555]=16'hfb1a;
aud[1556]=16'h9c81;
aud[1557]=16'h9962;
aud[1558]=16'hf49b;
aud[1559]=16'h5a4f;
aud[1560]=16'h6cfb;
aud[1561]=16'h1b75;
aud[1562]=16'hb0b1;
aud[1563]=16'h8ed7;
aud[1564]=16'hd508;
aud[1565]=16'h42ba;
aud[1566]=16'h7313;
aud[1567]=16'h39a0;
aud[1568]=16'hcb32;
aud[1569]=16'h8d51;
aud[1570]=16'hb8e0;
aud[1571]=16'h25d4;
aud[1572]=16'h7000;
aud[1573]=16'h5333;
aud[1574]=16'he9e8;
aud[1575]=16'h94ed;
aud[1576]=16'ha263;
aud[1577]=16'h5eb;
aud[1578]=16'h6402;
aud[1579]=16'h6626;
aud[1580]=16'ha61;
aud[1581]=16'ha510;
aud[1582]=16'h935b;
aud[1583]=16'he589;
aud[1584]=16'h500c;
aud[1585]=16'h70f6;
aud[1586]=16'h2a06;
aud[1587]=16'hbc72;
aud[1588]=16'h8cfb;
aud[1589]=16'hc743;
aud[1590]=16'h35b5;
aud[1591]=16'h72c7;
aud[1592]=16'h4652;
aud[1593]=16'hd936;
aud[1594]=16'h8fc4;
aud[1595]=16'had82;
aud[1596]=16'h1718;
aud[1597]=16'h6b72;
aud[1598]=16'h5d04;
aud[1599]=16'hf911;
aud[1600]=16'h9b7e;
aud[1601]=16'h9a53;
aud[1602]=16'hf6a3;
aud[1603]=16'h5b8f;
aud[1604]=16'h6c4d;
aud[1605]=16'h1979;
aud[1606]=16'haf39;
aud[1607]=16'h8f3e;
aud[1608]=16'hd6ee;
aud[1609]=16'h4460;
aud[1610]=16'h72f6;
aud[1611]=16'h37d9;
aud[1612]=16'hc964;
aud[1613]=16'h8d24;
aud[1614]=16'hba7e;
aud[1615]=16'h27bf;
aud[1616]=16'h7076;
aud[1617]=16'h51c7;
aud[1618]=16'he7e9;
aud[1619]=16'h9430;
aud[1620]=16'ha397;
aud[1621]=16'h7f4;
aud[1622]=16'h6501;
aud[1623]=16'h6531;
aud[1624]=16'h858;
aud[1625]=16'ha3d3;
aud[1626]=16'h940d;
aud[1627]=16'he786;
aud[1628]=16'h5180;
aud[1629]=16'h708c;
aud[1630]=16'h281e;
aud[1631]=16'hbace;
aud[1632]=16'h8d1c;
aud[1633]=16'hc90c;
aud[1634]=16'h3781;
aud[1635]=16'h72ef;
aud[1636]=16'h44b1;
aud[1637]=16'hd74c;
aud[1638]=16'h8f53;
aud[1639]=16'haef2;
aud[1640]=16'h1916;
aud[1641]=16'h6c2a;
aud[1642]=16'h5bcc;
aud[1643]=16'hf708;
aud[1644]=16'h9a83;
aud[1645]=16'h9b4d;
aud[1646]=16'hf8ac;
aud[1647]=16'h5cc8;
aud[1648]=16'h6b97;
aud[1649]=16'h177a;
aud[1650]=16'hadc8;
aud[1651]=16'h8fad;
aud[1652]=16'hd8d7;
aud[1653]=16'h4602;
aud[1654]=16'h72cf;
aud[1655]=16'h360e;
aud[1656]=16'hc79b;
aud[1657]=16'h8d01;
aud[1658]=16'hbc21;
aud[1659]=16'h29a8;
aud[1660]=16'h70e3;
aud[1661]=16'h5054;
aud[1662]=16'he5eb;
aud[1663]=16'h937d;
aud[1664]=16'ha4d3;
aud[1665]=16'h9fc;
aud[1666]=16'h65f8;
aud[1667]=16'h6433;
aud[1668]=16'h64f;
aud[1669]=16'ha29e;
aud[1670]=16'h94c8;
aud[1671]=16'he985;
aud[1672]=16'h52ee;
aud[1673]=16'h7018;
aud[1674]=16'h2633;
aud[1675]=16'hb930;
aud[1676]=16'h8d47;
aud[1677]=16'hcad9;
aud[1678]=16'h3948;
aud[1679]=16'h730e;
aud[1680]=16'h430b;
aud[1681]=16'hd565;
aud[1682]=16'h8eeb;
aud[1683]=16'hb068;
aud[1684]=16'h1b13;
aud[1685]=16'h6cda;
aud[1686]=16'h5a8d;
aud[1687]=16'hf500;
aud[1688]=16'h9990;
aud[1689]=16'h9c4e;
aud[1690]=16'hfab5;
aud[1691]=16'h5dfa;
aud[1692]=16'h6ad8;
aud[1693]=16'h157a;
aud[1694]=16'hac5e;
aud[1695]=16'h9026;
aud[1696]=16'hdac4;
aud[1697]=16'h479e;
aud[1698]=16'h72a0;
aud[1699]=16'h343f;
aud[1700]=16'hc5d6;
aud[1701]=16'h8ce6;
aud[1702]=16'hbdc9;
aud[1703]=16'h2b8d;
aud[1704]=16'h7146;
aud[1705]=16'h4edb;
aud[1706]=16'he3f0;
aud[1707]=16'h92d2;
aud[1708]=16'ha615;
aud[1709]=16'hc04;
aud[1710]=16'h66e7;
aud[1711]=16'h632e;
aud[1712]=16'h446;
aud[1713]=16'ha170;
aud[1714]=16'h958b;
aud[1715]=16'heb86;
aud[1716]=16'h5455;
aud[1717]=16'h6f9b;
aud[1718]=16'h2445;
aud[1719]=16'hb797;
aud[1720]=16'h8d7c;
aud[1721]=16'hccaa;
aud[1722]=16'h3b0b;
aud[1723]=16'h7323;
aud[1724]=16'h4160;
aud[1725]=16'hd382;
aud[1726]=16'h8e8b;
aud[1727]=16'hb1e5;
aud[1728]=16'h1d0d;
aud[1729]=16'h6d80;
aud[1730]=16'h5947;
aud[1731]=16'hf2f8;
aud[1732]=16'h98a5;
aud[1733]=16'h9d58;
aud[1734]=16'hfcbf;
aud[1735]=16'h5f24;
aud[1736]=16'h6a10;
aud[1737]=16'h1379;
aud[1738]=16'haafa;
aud[1739]=16'h90a7;
aud[1740]=16'hdcb3;
aud[1741]=16'h4934;
aud[1742]=16'h7267;
aud[1743]=16'h326c;
aud[1744]=16'hc415;
aud[1745]=16'h8cd5;
aud[1746]=16'hbf77;
aud[1747]=16'h2d6f;
aud[1748]=16'h71a1;
aud[1749]=16'h4d5b;
aud[1750]=16'he1f6;
aud[1751]=16'h9230;
aud[1752]=16'ha75f;
aud[1753]=16'he0b;
aud[1754]=16'h67cd;
aud[1755]=16'h6220;
aud[1756]=16'h23c;
aud[1757]=16'ha04a;
aud[1758]=16'h9657;
aud[1759]=16'hed89;
aud[1760]=16'h55b5;
aud[1761]=16'h6f15;
aud[1762]=16'h2254;
aud[1763]=16'hb603;
aud[1764]=16'h8db9;
aud[1765]=16'hce7f;
aud[1766]=16'h3cc9;
aud[1767]=16'h7330;
aud[1768]=16'h3fb0;
aud[1769]=16'hd1a2;
aud[1770]=16'h8e35;
aud[1771]=16'hb367;
aud[1772]=16'h1f05;
aud[1773]=16'h6e1e;
aud[1774]=16'h57f9;
aud[1775]=16'hf0f2;
aud[1776]=16'h97c3;
aud[1777]=16'h9e69;
aud[1778]=16'hfec9;
aud[1779]=16'h6047;
aud[1780]=16'h6940;
aud[1781]=16'h1175;
aud[1782]=16'ha99d;
aud[1783]=16'h9132;
aud[1784]=16'hdea6;
aud[1785]=16'h4ac4;
aud[1786]=16'h7225;
aud[1787]=16'h3094;
aud[1788]=16'hc25a;
aud[1789]=16'h8ccd;
aud[1790]=16'hc12a;
aud[1791]=16'h2f4c;
aud[1792]=16'h71f2;
aud[1793]=16'h4bd5;
aud[1794]=16'he000;
aud[1795]=16'h9196;
aud[1796]=16'ha8b0;
aud[1797]=16'h1010;
aud[1798]=16'h68ab;
aud[1799]=16'h610b;
aud[1800]=16'h32;
aud[1801]=16'h9f2b;
aud[1802]=16'h972b;
aud[1803]=16'hef8d;
aud[1804]=16'h570e;
aud[1805]=16'h6e86;
aud[1806]=16'h2060;
aud[1807]=16'hb476;
aud[1808]=16'h8dff;
aud[1809]=16'hd059;
aud[1810]=16'h3e82;
aud[1811]=16'h7333;
aud[1812]=16'h3dfa;
aud[1813]=16'hcfc6;
aud[1814]=16'h8de9;
aud[1815]=16'hb4f0;
aud[1816]=16'h20fb;
aud[1817]=16'h6eb3;
aud[1818]=16'h56a4;
aud[1819]=16'heeed;
aud[1820]=16'h96e9;
aud[1821]=16'h9f83;
aud[1822]=16'hd3;
aud[1823]=16'h6161;
aud[1824]=16'h6868;
aud[1825]=16'hf71;
aud[1826]=16'ha848;
aud[1827]=16'h91c5;
aud[1828]=16'he09b;
aud[1829]=16'h4c4e;
aud[1830]=16'h71da;
aud[1831]=16'h2eb9;
aud[1832]=16'hc0a3;
aud[1833]=16'h8ccf;
aud[1834]=16'hc2e2;
aud[1835]=16'h3127;
aud[1836]=16'h723a;
aud[1837]=16'h4a49;
aud[1838]=16'hde0b;
aud[1839]=16'h9106;
aud[1840]=16'haa08;
aud[1841]=16'h1215;
aud[1842]=16'h6981;
aud[1843]=16'h5fee;
aud[1844]=16'hfe28;
aud[1845]=16'h9e14;
aud[1846]=16'h9808;
aud[1847]=16'hf192;
aud[1848]=16'h5861;
aud[1849]=16'h6dee;
aud[1850]=16'h1e6a;
aud[1851]=16'hb2ef;
aud[1852]=16'h8e4f;
aud[1853]=16'hd236;
aud[1854]=16'h4036;
aud[1855]=16'h732d;
aud[1856]=16'h3c40;
aud[1857]=16'hcdee;
aud[1858]=16'h8da5;
aud[1859]=16'hb67f;
aud[1860]=16'h22ee;
aud[1861]=16'h6f3f;
aud[1862]=16'h5549;
aud[1863]=16'hecea;
aud[1864]=16'h9617;
aud[1865]=16'ha0a4;
aud[1866]=16'h2dd;
aud[1867]=16'h6274;
aud[1868]=16'h6787;
aud[1869]=16'hd6b;
aud[1870]=16'ha6f9;
aud[1871]=16'h9261;
aud[1872]=16'he292;
aud[1873]=16'h4dd2;
aud[1874]=16'h7186;
aud[1875]=16'h2cda;
aud[1876]=16'hbef2;
aud[1877]=16'h8cd9;
aud[1878]=16'hc49f;
aud[1879]=16'h32fd;
aud[1880]=16'h7279;
aud[1881]=16'h48b7;
aud[1882]=16'hdc1a;
aud[1883]=16'h907e;
aud[1884]=16'hab67;
aud[1885]=16'h1418;
aud[1886]=16'h6a4f;
aud[1887]=16'h5ec9;
aud[1888]=16'hfc1e;
aud[1889]=16'h9d05;
aud[1890]=16'h98ed;
aud[1891]=16'hf399;
aud[1892]=16'h59ac;
aud[1893]=16'h6d4e;
aud[1894]=16'h1c71;
aud[1895]=16'hb16e;
aud[1896]=16'h8ea8;
aud[1897]=16'hd417;
aud[1898]=16'h41e5;
aud[1899]=16'h731e;
aud[1900]=16'h3a80;
aud[1901]=16'hcc1a;
aud[1902]=16'h8d6a;
aud[1903]=16'hb814;
aud[1904]=16'h24de;
aud[1905]=16'h6fc2;
aud[1906]=16'h53e7;
aud[1907]=16'heae8;
aud[1908]=16'h954e;
aud[1909]=16'ha1cd;
aud[1910]=16'h4e7;
aud[1911]=16'h6380;
aud[1912]=16'h669e;
aud[1913]=16'hb64;
aud[1914]=16'ha5b1;
aud[1915]=16'h9306;
aud[1916]=16'he48c;
aud[1917]=16'h4f50;
aud[1918]=16'h7128;
aud[1919]=16'h2af7;
aud[1920]=16'hbd46;
aud[1921]=16'h8ced;
aud[1922]=16'hc661;
aud[1923]=16'h34cf;
aud[1924]=16'h72af;
aud[1925]=16'h471f;
aud[1926]=16'hda2b;
aud[1927]=16'h9000;
aud[1928]=16'haccd;
aud[1929]=16'h1619;
aud[1930]=16'h6b14;
aud[1931]=16'h5d9c;
aud[1932]=16'hfa14;
aud[1933]=16'h9bfe;
aud[1934]=16'h99da;
aud[1935]=16'hf5a0;
aud[1936]=16'h5af0;
aud[1937]=16'h6ca5;
aud[1938]=16'h1a76;
aud[1939]=16'haff4;
aud[1940]=16'h8f0a;
aud[1941]=16'hd5fb;
aud[1942]=16'h438e;
aud[1943]=16'h7305;
aud[1944]=16'h38bc;
aud[1945]=16'hca4a;
aud[1946]=16'h8d39;
aud[1947]=16'hb9af;
aud[1948]=16'h26cb;
aud[1949]=16'h703c;
aud[1950]=16'h527d;
aud[1951]=16'he8e7;
aud[1952]=16'h948d;
aud[1953]=16'ha2fd;
aud[1954]=16'h6f0;
aud[1955]=16'h6483;
aud[1956]=16'h65ac;
aud[1957]=16'h95c;
aud[1958]=16'ha470;
aud[1959]=16'h93b3;
aud[1960]=16'he688;
aud[1961]=16'h50c7;
aud[1962]=16'h70c2;
aud[1963]=16'h2911;
aud[1964]=16'hbb9f;
aud[1965]=16'h8d0a;
aud[1966]=16'hc828;
aud[1967]=16'h369d;
aud[1968]=16'h72dc;
aud[1969]=16'h4581;
aud[1970]=16'hd840;
aud[1971]=16'h8f8a;
aud[1972]=16'hae3a;
aud[1973]=16'h1818;
aud[1974]=16'h6bd0;
aud[1975]=16'h5c68;
aud[1976]=16'hf80b;
aud[1977]=16'h9aff;
aud[1978]=16'h9acf;
aud[1979]=16'hf7a9;
aud[1980]=16'h5c2d;
aud[1981]=16'h6bf3;
aud[1982]=16'h1879;
aud[1983]=16'hae7f;
aud[1984]=16'h8f75;
aud[1985]=16'hd7e3;
aud[1986]=16'h4533;
aud[1987]=16'h72e3;
aud[1988]=16'h36f4;
aud[1989]=16'hc87e;
aud[1990]=16'h8d11;
aud[1991]=16'hbb4f;
aud[1992]=16'h28b5;
aud[1993]=16'h70ae;
aud[1994]=16'h510e;
aud[1995]=16'he6e9;
aud[1996]=16'h93d5;
aud[1997]=16'ha435;
aud[1998]=16'h8f9;
aud[1999]=16'h657e;

end


endmodule