module testVect (
output reg signed [15:0] aud [0:1999]
);

initial begin
aud[0]=16'hf09;
aud[1]=16'h1dd1;
aud[2]=16'h2c16;
aud[3]=16'h399a;
aud[4]=16'h4621;
aud[5]=16'h5175;
aud[6]=16'h5b65;
aud[7]=16'h63c4;
aud[8]=16'h6a6e;
aud[9]=16'h6f46;
aud[10]=16'h7237;
aud[11]=16'h7333;
aud[12]=16'h7237;
aud[13]=16'h6f46;
aud[14]=16'h6a6e;
aud[15]=16'h63c4;
aud[16]=16'h5b65;
aud[17]=16'h5175;
aud[18]=16'h4621;
aud[19]=16'h399a;
aud[20]=16'h2c16;
aud[21]=16'h1dd1;
aud[22]=16'hf09;
aud[23]=16'h0;
aud[24]=16'hf0f7;
aud[25]=16'he22f;
aud[26]=16'hd3ea;
aud[27]=16'hc666;
aud[28]=16'hb9df;
aud[29]=16'hae8b;
aud[30]=16'ha49b;
aud[31]=16'h9c3c;
aud[32]=16'h9592;
aud[33]=16'h90ba;
aud[34]=16'h8dc9;
aud[35]=16'h8ccd;
aud[36]=16'h8dc9;
aud[37]=16'h90ba;
aud[38]=16'h9592;
aud[39]=16'h9c3c;
aud[40]=16'ha49b;
aud[41]=16'hae8b;
aud[42]=16'hb9df;
aud[43]=16'hc666;
aud[44]=16'hd3ea;
aud[45]=16'he22f;
aud[46]=16'hf0f7;
aud[47]=16'h0;
aud[48]=16'hf09;
aud[49]=16'h1dd1;
aud[50]=16'h2c16;
aud[51]=16'h399a;
aud[52]=16'h4621;
aud[53]=16'h5175;
aud[54]=16'h5b65;
aud[55]=16'h63c4;
aud[56]=16'h6a6e;
aud[57]=16'h6f46;
aud[58]=16'h7237;
aud[59]=16'h7333;
aud[60]=16'h7237;
aud[61]=16'h6f46;
aud[62]=16'h6a6e;
aud[63]=16'h63c4;
aud[64]=16'h5b65;
aud[65]=16'h5175;
aud[66]=16'h4621;
aud[67]=16'h399a;
aud[68]=16'h2c16;
aud[69]=16'h1dd1;
aud[70]=16'hf09;
aud[71]=16'h0;
aud[72]=16'hf0f7;
aud[73]=16'he22f;
aud[74]=16'hd3ea;
aud[75]=16'hc666;
aud[76]=16'hb9df;
aud[77]=16'hae8b;
aud[78]=16'ha49b;
aud[79]=16'h9c3c;
aud[80]=16'h9592;
aud[81]=16'h90ba;
aud[82]=16'h8dc9;
aud[83]=16'h8ccd;
aud[84]=16'h8dc9;
aud[85]=16'h90ba;
aud[86]=16'h9592;
aud[87]=16'h9c3c;
aud[88]=16'ha49b;
aud[89]=16'hae8b;
aud[90]=16'hb9df;
aud[91]=16'hc666;
aud[92]=16'hd3ea;
aud[93]=16'he22f;
aud[94]=16'hf0f7;
aud[95]=16'h0;
aud[96]=16'hf09;
aud[97]=16'h1dd1;
aud[98]=16'h2c16;
aud[99]=16'h399a;
aud[100]=16'h4621;
aud[101]=16'h5175;
aud[102]=16'h5b65;
aud[103]=16'h63c4;
aud[104]=16'h6a6e;
aud[105]=16'h6f46;
aud[106]=16'h7237;
aud[107]=16'h7333;
aud[108]=16'h7237;
aud[109]=16'h6f46;
aud[110]=16'h6a6e;
aud[111]=16'h63c4;
aud[112]=16'h5b65;
aud[113]=16'h5175;
aud[114]=16'h4621;
aud[115]=16'h399a;
aud[116]=16'h2c16;
aud[117]=16'h1dd1;
aud[118]=16'hf09;
aud[119]=16'h0;
aud[120]=16'hf0f7;
aud[121]=16'he22f;
aud[122]=16'hd3ea;
aud[123]=16'hc666;
aud[124]=16'hb9df;
aud[125]=16'hae8b;
aud[126]=16'ha49b;
aud[127]=16'h9c3c;
aud[128]=16'h9592;
aud[129]=16'h90ba;
aud[130]=16'h8dc9;
aud[131]=16'h8ccd;
aud[132]=16'h8dc9;
aud[133]=16'h90ba;
aud[134]=16'h9592;
aud[135]=16'h9c3c;
aud[136]=16'ha49b;
aud[137]=16'hae8b;
aud[138]=16'hb9df;
aud[139]=16'hc666;
aud[140]=16'hd3ea;
aud[141]=16'he22f;
aud[142]=16'hf0f7;
aud[143]=16'h0;
aud[144]=16'hf09;
aud[145]=16'h1dd1;
aud[146]=16'h2c16;
aud[147]=16'h399a;
aud[148]=16'h4621;
aud[149]=16'h5175;
aud[150]=16'h5b65;
aud[151]=16'h63c4;
aud[152]=16'h6a6e;
aud[153]=16'h6f46;
aud[154]=16'h7237;
aud[155]=16'h7333;
aud[156]=16'h7237;
aud[157]=16'h6f46;
aud[158]=16'h6a6e;
aud[159]=16'h63c4;
aud[160]=16'h5b65;
aud[161]=16'h5175;
aud[162]=16'h4621;
aud[163]=16'h399a;
aud[164]=16'h2c16;
aud[165]=16'h1dd1;
aud[166]=16'hf09;
aud[167]=16'h0;
aud[168]=16'hf0f7;
aud[169]=16'he22f;
aud[170]=16'hd3ea;
aud[171]=16'hc666;
aud[172]=16'hb9df;
aud[173]=16'hae8b;
aud[174]=16'ha49b;
aud[175]=16'h9c3c;
aud[176]=16'h9592;
aud[177]=16'h90ba;
aud[178]=16'h8dc9;
aud[179]=16'h8ccd;
aud[180]=16'h8dc9;
aud[181]=16'h90ba;
aud[182]=16'h9592;
aud[183]=16'h9c3c;
aud[184]=16'ha49b;
aud[185]=16'hae8b;
aud[186]=16'hb9df;
aud[187]=16'hc666;
aud[188]=16'hd3ea;
aud[189]=16'he22f;
aud[190]=16'hf0f7;
aud[191]=16'h0;
aud[192]=16'hf09;
aud[193]=16'h1dd1;
aud[194]=16'h2c16;
aud[195]=16'h399a;
aud[196]=16'h4621;
aud[197]=16'h5175;
aud[198]=16'h5b65;
aud[199]=16'h63c4;
aud[200]=16'h6a6e;
aud[201]=16'h6f46;
aud[202]=16'h7237;
aud[203]=16'h7333;
aud[204]=16'h7237;
aud[205]=16'h6f46;
aud[206]=16'h6a6e;
aud[207]=16'h63c4;
aud[208]=16'h5b65;
aud[209]=16'h5175;
aud[210]=16'h4621;
aud[211]=16'h399a;
aud[212]=16'h2c16;
aud[213]=16'h1dd1;
aud[214]=16'hf09;
aud[215]=16'h0;
aud[216]=16'hf0f7;
aud[217]=16'he22f;
aud[218]=16'hd3ea;
aud[219]=16'hc666;
aud[220]=16'hb9df;
aud[221]=16'hae8b;
aud[222]=16'ha49b;
aud[223]=16'h9c3c;
aud[224]=16'h9592;
aud[225]=16'h90ba;
aud[226]=16'h8dc9;
aud[227]=16'h8ccd;
aud[228]=16'h8dc9;
aud[229]=16'h90ba;
aud[230]=16'h9592;
aud[231]=16'h9c3c;
aud[232]=16'ha49b;
aud[233]=16'hae8b;
aud[234]=16'hb9df;
aud[235]=16'hc666;
aud[236]=16'hd3ea;
aud[237]=16'he22f;
aud[238]=16'hf0f7;
aud[239]=16'h0;
aud[240]=16'hf09;
aud[241]=16'h1dd1;
aud[242]=16'h2c16;
aud[243]=16'h399a;
aud[244]=16'h4621;
aud[245]=16'h5175;
aud[246]=16'h5b65;
aud[247]=16'h63c4;
aud[248]=16'h6a6e;
aud[249]=16'h6f46;
aud[250]=16'h7237;
aud[251]=16'h7333;
aud[252]=16'h7237;
aud[253]=16'h6f46;
aud[254]=16'h6a6e;
aud[255]=16'h63c4;
aud[256]=16'h5b65;
aud[257]=16'h5175;
aud[258]=16'h4621;
aud[259]=16'h399a;
aud[260]=16'h2c16;
aud[261]=16'h1dd1;
aud[262]=16'hf09;
aud[263]=16'h0;
aud[264]=16'hf0f7;
aud[265]=16'he22f;
aud[266]=16'hd3ea;
aud[267]=16'hc666;
aud[268]=16'hb9df;
aud[269]=16'hae8b;
aud[270]=16'ha49b;
aud[271]=16'h9c3c;
aud[272]=16'h9592;
aud[273]=16'h90ba;
aud[274]=16'h8dc9;
aud[275]=16'h8ccd;
aud[276]=16'h8dc9;
aud[277]=16'h90ba;
aud[278]=16'h9592;
aud[279]=16'h9c3c;
aud[280]=16'ha49b;
aud[281]=16'hae8b;
aud[282]=16'hb9df;
aud[283]=16'hc666;
aud[284]=16'hd3ea;
aud[285]=16'he22f;
aud[286]=16'hf0f7;
aud[287]=16'h0;
aud[288]=16'hf09;
aud[289]=16'h1dd1;
aud[290]=16'h2c16;
aud[291]=16'h399a;
aud[292]=16'h4621;
aud[293]=16'h5175;
aud[294]=16'h5b65;
aud[295]=16'h63c4;
aud[296]=16'h6a6e;
aud[297]=16'h6f46;
aud[298]=16'h7237;
aud[299]=16'h7333;
aud[300]=16'h7237;
aud[301]=16'h6f46;
aud[302]=16'h6a6e;
aud[303]=16'h63c4;
aud[304]=16'h5b65;
aud[305]=16'h5175;
aud[306]=16'h4621;
aud[307]=16'h399a;
aud[308]=16'h2c16;
aud[309]=16'h1dd1;
aud[310]=16'hf09;
aud[311]=16'h0;
aud[312]=16'hf0f7;
aud[313]=16'he22f;
aud[314]=16'hd3ea;
aud[315]=16'hc666;
aud[316]=16'hb9df;
aud[317]=16'hae8b;
aud[318]=16'ha49b;
aud[319]=16'h9c3c;
aud[320]=16'h9592;
aud[321]=16'h90ba;
aud[322]=16'h8dc9;
aud[323]=16'h8ccd;
aud[324]=16'h8dc9;
aud[325]=16'h90ba;
aud[326]=16'h9592;
aud[327]=16'h9c3c;
aud[328]=16'ha49b;
aud[329]=16'hae8b;
aud[330]=16'hb9df;
aud[331]=16'hc666;
aud[332]=16'hd3ea;
aud[333]=16'he22f;
aud[334]=16'hf0f7;
aud[335]=16'h0;
aud[336]=16'hf09;
aud[337]=16'h1dd1;
aud[338]=16'h2c16;
aud[339]=16'h399a;
aud[340]=16'h4621;
aud[341]=16'h5175;
aud[342]=16'h5b65;
aud[343]=16'h63c4;
aud[344]=16'h6a6e;
aud[345]=16'h6f46;
aud[346]=16'h7237;
aud[347]=16'h7333;
aud[348]=16'h7237;
aud[349]=16'h6f46;
aud[350]=16'h6a6e;
aud[351]=16'h63c4;
aud[352]=16'h5b65;
aud[353]=16'h5175;
aud[354]=16'h4621;
aud[355]=16'h399a;
aud[356]=16'h2c16;
aud[357]=16'h1dd1;
aud[358]=16'hf09;
aud[359]=16'h0;
aud[360]=16'hf0f7;
aud[361]=16'he22f;
aud[362]=16'hd3ea;
aud[363]=16'hc666;
aud[364]=16'hb9df;
aud[365]=16'hae8b;
aud[366]=16'ha49b;
aud[367]=16'h9c3c;
aud[368]=16'h9592;
aud[369]=16'h90ba;
aud[370]=16'h8dc9;
aud[371]=16'h8ccd;
aud[372]=16'h8dc9;
aud[373]=16'h90ba;
aud[374]=16'h9592;
aud[375]=16'h9c3c;
aud[376]=16'ha49b;
aud[377]=16'hae8b;
aud[378]=16'hb9df;
aud[379]=16'hc666;
aud[380]=16'hd3ea;
aud[381]=16'he22f;
aud[382]=16'hf0f7;
aud[383]=16'h0;
aud[384]=16'hf09;
aud[385]=16'h1dd1;
aud[386]=16'h2c16;
aud[387]=16'h399a;
aud[388]=16'h4621;
aud[389]=16'h5175;
aud[390]=16'h5b65;
aud[391]=16'h63c4;
aud[392]=16'h6a6e;
aud[393]=16'h6f46;
aud[394]=16'h7237;
aud[395]=16'h7333;
aud[396]=16'h7237;
aud[397]=16'h6f46;
aud[398]=16'h6a6e;
aud[399]=16'h63c4;
aud[400]=16'h5b65;
aud[401]=16'h5175;
aud[402]=16'h4621;
aud[403]=16'h399a;
aud[404]=16'h2c16;
aud[405]=16'h1dd1;
aud[406]=16'hf09;
aud[407]=16'h0;
aud[408]=16'hf0f7;
aud[409]=16'he22f;
aud[410]=16'hd3ea;
aud[411]=16'hc666;
aud[412]=16'hb9df;
aud[413]=16'hae8b;
aud[414]=16'ha49b;
aud[415]=16'h9c3c;
aud[416]=16'h9592;
aud[417]=16'h90ba;
aud[418]=16'h8dc9;
aud[419]=16'h8ccd;
aud[420]=16'h8dc9;
aud[421]=16'h90ba;
aud[422]=16'h9592;
aud[423]=16'h9c3c;
aud[424]=16'ha49b;
aud[425]=16'hae8b;
aud[426]=16'hb9df;
aud[427]=16'hc666;
aud[428]=16'hd3ea;
aud[429]=16'he22f;
aud[430]=16'hf0f7;
aud[431]=16'h0;
aud[432]=16'hf09;
aud[433]=16'h1dd1;
aud[434]=16'h2c16;
aud[435]=16'h399a;
aud[436]=16'h4621;
aud[437]=16'h5175;
aud[438]=16'h5b65;
aud[439]=16'h63c4;
aud[440]=16'h6a6e;
aud[441]=16'h6f46;
aud[442]=16'h7237;
aud[443]=16'h7333;
aud[444]=16'h7237;
aud[445]=16'h6f46;
aud[446]=16'h6a6e;
aud[447]=16'h63c4;
aud[448]=16'h5b65;
aud[449]=16'h5175;
aud[450]=16'h4621;
aud[451]=16'h399a;
aud[452]=16'h2c16;
aud[453]=16'h1dd1;
aud[454]=16'hf09;
aud[455]=16'h0;
aud[456]=16'hf0f7;
aud[457]=16'he22f;
aud[458]=16'hd3ea;
aud[459]=16'hc666;
aud[460]=16'hb9df;
aud[461]=16'hae8b;
aud[462]=16'ha49b;
aud[463]=16'h9c3c;
aud[464]=16'h9592;
aud[465]=16'h90ba;
aud[466]=16'h8dc9;
aud[467]=16'h8ccd;
aud[468]=16'h8dc9;
aud[469]=16'h90ba;
aud[470]=16'h9592;
aud[471]=16'h9c3c;
aud[472]=16'ha49b;
aud[473]=16'hae8b;
aud[474]=16'hb9df;
aud[475]=16'hc666;
aud[476]=16'hd3ea;
aud[477]=16'he22f;
aud[478]=16'hf0f7;
aud[479]=16'h0;
aud[480]=16'hf09;
aud[481]=16'h1dd1;
aud[482]=16'h2c16;
aud[483]=16'h399a;
aud[484]=16'h4621;
aud[485]=16'h5175;
aud[486]=16'h5b65;
aud[487]=16'h63c4;
aud[488]=16'h6a6e;
aud[489]=16'h6f46;
aud[490]=16'h7237;
aud[491]=16'h7333;
aud[492]=16'h7237;
aud[493]=16'h6f46;
aud[494]=16'h6a6e;
aud[495]=16'h63c4;
aud[496]=16'h5b65;
aud[497]=16'h5175;
aud[498]=16'h4621;
aud[499]=16'h399a;
aud[500]=16'h2c16;
aud[501]=16'h1dd1;
aud[502]=16'hf09;
aud[503]=16'h0;
aud[504]=16'hf0f7;
aud[505]=16'he22f;
aud[506]=16'hd3ea;
aud[507]=16'hc666;
aud[508]=16'hb9df;
aud[509]=16'hae8b;
aud[510]=16'ha49b;
aud[511]=16'h9c3c;
aud[512]=16'h9592;
aud[513]=16'h90ba;
aud[514]=16'h8dc9;
aud[515]=16'h8ccd;
aud[516]=16'h8dc9;
aud[517]=16'h90ba;
aud[518]=16'h9592;
aud[519]=16'h9c3c;
aud[520]=16'ha49b;
aud[521]=16'hae8b;
aud[522]=16'hb9df;
aud[523]=16'hc666;
aud[524]=16'hd3ea;
aud[525]=16'he22f;
aud[526]=16'hf0f7;
aud[527]=16'h0;
aud[528]=16'hf09;
aud[529]=16'h1dd1;
aud[530]=16'h2c16;
aud[531]=16'h399a;
aud[532]=16'h4621;
aud[533]=16'h5175;
aud[534]=16'h5b65;
aud[535]=16'h63c4;
aud[536]=16'h6a6e;
aud[537]=16'h6f46;
aud[538]=16'h7237;
aud[539]=16'h7333;
aud[540]=16'h7237;
aud[541]=16'h6f46;
aud[542]=16'h6a6e;
aud[543]=16'h63c4;
aud[544]=16'h5b65;
aud[545]=16'h5175;
aud[546]=16'h4621;
aud[547]=16'h399a;
aud[548]=16'h2c16;
aud[549]=16'h1dd1;
aud[550]=16'hf09;
aud[551]=16'h0;
aud[552]=16'hf0f7;
aud[553]=16'he22f;
aud[554]=16'hd3ea;
aud[555]=16'hc666;
aud[556]=16'hb9df;
aud[557]=16'hae8b;
aud[558]=16'ha49b;
aud[559]=16'h9c3c;
aud[560]=16'h9592;
aud[561]=16'h90ba;
aud[562]=16'h8dc9;
aud[563]=16'h8ccd;
aud[564]=16'h8dc9;
aud[565]=16'h90ba;
aud[566]=16'h9592;
aud[567]=16'h9c3c;
aud[568]=16'ha49b;
aud[569]=16'hae8b;
aud[570]=16'hb9df;
aud[571]=16'hc666;
aud[572]=16'hd3ea;
aud[573]=16'he22f;
aud[574]=16'hf0f7;
aud[575]=16'h0;
aud[576]=16'hf09;
aud[577]=16'h1dd1;
aud[578]=16'h2c16;
aud[579]=16'h399a;
aud[580]=16'h4621;
aud[581]=16'h5175;
aud[582]=16'h5b65;
aud[583]=16'h63c4;
aud[584]=16'h6a6e;
aud[585]=16'h6f46;
aud[586]=16'h7237;
aud[587]=16'h7333;
aud[588]=16'h7237;
aud[589]=16'h6f46;
aud[590]=16'h6a6e;
aud[591]=16'h63c4;
aud[592]=16'h5b65;
aud[593]=16'h5175;
aud[594]=16'h4621;
aud[595]=16'h399a;
aud[596]=16'h2c16;
aud[597]=16'h1dd1;
aud[598]=16'hf09;
aud[599]=16'h0;
aud[600]=16'hf0f7;
aud[601]=16'he22f;
aud[602]=16'hd3ea;
aud[603]=16'hc666;
aud[604]=16'hb9df;
aud[605]=16'hae8b;
aud[606]=16'ha49b;
aud[607]=16'h9c3c;
aud[608]=16'h9592;
aud[609]=16'h90ba;
aud[610]=16'h8dc9;
aud[611]=16'h8ccd;
aud[612]=16'h8dc9;
aud[613]=16'h90ba;
aud[614]=16'h9592;
aud[615]=16'h9c3c;
aud[616]=16'ha49b;
aud[617]=16'hae8b;
aud[618]=16'hb9df;
aud[619]=16'hc666;
aud[620]=16'hd3ea;
aud[621]=16'he22f;
aud[622]=16'hf0f7;
aud[623]=16'h0;
aud[624]=16'hf09;
aud[625]=16'h1dd1;
aud[626]=16'h2c16;
aud[627]=16'h399a;
aud[628]=16'h4621;
aud[629]=16'h5175;
aud[630]=16'h5b65;
aud[631]=16'h63c4;
aud[632]=16'h6a6e;
aud[633]=16'h6f46;
aud[634]=16'h7237;
aud[635]=16'h7333;
aud[636]=16'h7237;
aud[637]=16'h6f46;
aud[638]=16'h6a6e;
aud[639]=16'h63c4;
aud[640]=16'h5b65;
aud[641]=16'h5175;
aud[642]=16'h4621;
aud[643]=16'h399a;
aud[644]=16'h2c16;
aud[645]=16'h1dd1;
aud[646]=16'hf09;
aud[647]=16'h0;
aud[648]=16'hf0f7;
aud[649]=16'he22f;
aud[650]=16'hd3ea;
aud[651]=16'hc666;
aud[652]=16'hb9df;
aud[653]=16'hae8b;
aud[654]=16'ha49b;
aud[655]=16'h9c3c;
aud[656]=16'h9592;
aud[657]=16'h90ba;
aud[658]=16'h8dc9;
aud[659]=16'h8ccd;
aud[660]=16'h8dc9;
aud[661]=16'h90ba;
aud[662]=16'h9592;
aud[663]=16'h9c3c;
aud[664]=16'ha49b;
aud[665]=16'hae8b;
aud[666]=16'hb9df;
aud[667]=16'hc666;
aud[668]=16'hd3ea;
aud[669]=16'he22f;
aud[670]=16'hf0f7;
aud[671]=16'h0;
aud[672]=16'hf09;
aud[673]=16'h1dd1;
aud[674]=16'h2c16;
aud[675]=16'h399a;
aud[676]=16'h4621;
aud[677]=16'h5175;
aud[678]=16'h5b65;
aud[679]=16'h63c4;
aud[680]=16'h6a6e;
aud[681]=16'h6f46;
aud[682]=16'h7237;
aud[683]=16'h7333;
aud[684]=16'h7237;
aud[685]=16'h6f46;
aud[686]=16'h6a6e;
aud[687]=16'h63c4;
aud[688]=16'h5b65;
aud[689]=16'h5175;
aud[690]=16'h4621;
aud[691]=16'h399a;
aud[692]=16'h2c16;
aud[693]=16'h1dd1;
aud[694]=16'hf09;
aud[695]=16'h0;
aud[696]=16'hf0f7;
aud[697]=16'he22f;
aud[698]=16'hd3ea;
aud[699]=16'hc666;
aud[700]=16'hb9df;
aud[701]=16'hae8b;
aud[702]=16'ha49b;
aud[703]=16'h9c3c;
aud[704]=16'h9592;
aud[705]=16'h90ba;
aud[706]=16'h8dc9;
aud[707]=16'h8ccd;
aud[708]=16'h8dc9;
aud[709]=16'h90ba;
aud[710]=16'h9592;
aud[711]=16'h9c3c;
aud[712]=16'ha49b;
aud[713]=16'hae8b;
aud[714]=16'hb9df;
aud[715]=16'hc666;
aud[716]=16'hd3ea;
aud[717]=16'he22f;
aud[718]=16'hf0f7;
aud[719]=16'h0;
aud[720]=16'hf09;
aud[721]=16'h1dd1;
aud[722]=16'h2c16;
aud[723]=16'h399a;
aud[724]=16'h4621;
aud[725]=16'h5175;
aud[726]=16'h5b65;
aud[727]=16'h63c4;
aud[728]=16'h6a6e;
aud[729]=16'h6f46;
aud[730]=16'h7237;
aud[731]=16'h7333;
aud[732]=16'h7237;
aud[733]=16'h6f46;
aud[734]=16'h6a6e;
aud[735]=16'h63c4;
aud[736]=16'h5b65;
aud[737]=16'h5175;
aud[738]=16'h4621;
aud[739]=16'h399a;
aud[740]=16'h2c16;
aud[741]=16'h1dd1;
aud[742]=16'hf09;
aud[743]=16'h0;
aud[744]=16'hf0f7;
aud[745]=16'he22f;
aud[746]=16'hd3ea;
aud[747]=16'hc666;
aud[748]=16'hb9df;
aud[749]=16'hae8b;
aud[750]=16'ha49b;
aud[751]=16'h9c3c;
aud[752]=16'h9592;
aud[753]=16'h90ba;
aud[754]=16'h8dc9;
aud[755]=16'h8ccd;
aud[756]=16'h8dc9;
aud[757]=16'h90ba;
aud[758]=16'h9592;
aud[759]=16'h9c3c;
aud[760]=16'ha49b;
aud[761]=16'hae8b;
aud[762]=16'hb9df;
aud[763]=16'hc666;
aud[764]=16'hd3ea;
aud[765]=16'he22f;
aud[766]=16'hf0f7;
aud[767]=16'h0;
aud[768]=16'hf09;
aud[769]=16'h1dd1;
aud[770]=16'h2c16;
aud[771]=16'h399a;
aud[772]=16'h4621;
aud[773]=16'h5175;
aud[774]=16'h5b65;
aud[775]=16'h63c4;
aud[776]=16'h6a6e;
aud[777]=16'h6f46;
aud[778]=16'h7237;
aud[779]=16'h7333;
aud[780]=16'h7237;
aud[781]=16'h6f46;
aud[782]=16'h6a6e;
aud[783]=16'h63c4;
aud[784]=16'h5b65;
aud[785]=16'h5175;
aud[786]=16'h4621;
aud[787]=16'h399a;
aud[788]=16'h2c16;
aud[789]=16'h1dd1;
aud[790]=16'hf09;
aud[791]=16'h0;
aud[792]=16'hf0f7;
aud[793]=16'he22f;
aud[794]=16'hd3ea;
aud[795]=16'hc666;
aud[796]=16'hb9df;
aud[797]=16'hae8b;
aud[798]=16'ha49b;
aud[799]=16'h9c3c;
aud[800]=16'h9592;
aud[801]=16'h90ba;
aud[802]=16'h8dc9;
aud[803]=16'h8ccd;
aud[804]=16'h8dc9;
aud[805]=16'h90ba;
aud[806]=16'h9592;
aud[807]=16'h9c3c;
aud[808]=16'ha49b;
aud[809]=16'hae8b;
aud[810]=16'hb9df;
aud[811]=16'hc666;
aud[812]=16'hd3ea;
aud[813]=16'he22f;
aud[814]=16'hf0f7;
aud[815]=16'h0;
aud[816]=16'hf09;
aud[817]=16'h1dd1;
aud[818]=16'h2c16;
aud[819]=16'h399a;
aud[820]=16'h4621;
aud[821]=16'h5175;
aud[822]=16'h5b65;
aud[823]=16'h63c4;
aud[824]=16'h6a6e;
aud[825]=16'h6f46;
aud[826]=16'h7237;
aud[827]=16'h7333;
aud[828]=16'h7237;
aud[829]=16'h6f46;
aud[830]=16'h6a6e;
aud[831]=16'h63c4;
aud[832]=16'h5b65;
aud[833]=16'h5175;
aud[834]=16'h4621;
aud[835]=16'h399a;
aud[836]=16'h2c16;
aud[837]=16'h1dd1;
aud[838]=16'hf09;
aud[839]=16'h0;
aud[840]=16'hf0f7;
aud[841]=16'he22f;
aud[842]=16'hd3ea;
aud[843]=16'hc666;
aud[844]=16'hb9df;
aud[845]=16'hae8b;
aud[846]=16'ha49b;
aud[847]=16'h9c3c;
aud[848]=16'h9592;
aud[849]=16'h90ba;
aud[850]=16'h8dc9;
aud[851]=16'h8ccd;
aud[852]=16'h8dc9;
aud[853]=16'h90ba;
aud[854]=16'h9592;
aud[855]=16'h9c3c;
aud[856]=16'ha49b;
aud[857]=16'hae8b;
aud[858]=16'hb9df;
aud[859]=16'hc666;
aud[860]=16'hd3ea;
aud[861]=16'he22f;
aud[862]=16'hf0f7;
aud[863]=16'h0;
aud[864]=16'hf09;
aud[865]=16'h1dd1;
aud[866]=16'h2c16;
aud[867]=16'h399a;
aud[868]=16'h4621;
aud[869]=16'h5175;
aud[870]=16'h5b65;
aud[871]=16'h63c4;
aud[872]=16'h6a6e;
aud[873]=16'h6f46;
aud[874]=16'h7237;
aud[875]=16'h7333;
aud[876]=16'h7237;
aud[877]=16'h6f46;
aud[878]=16'h6a6e;
aud[879]=16'h63c4;
aud[880]=16'h5b65;
aud[881]=16'h5175;
aud[882]=16'h4621;
aud[883]=16'h399a;
aud[884]=16'h2c16;
aud[885]=16'h1dd1;
aud[886]=16'hf09;
aud[887]=16'h0;
aud[888]=16'hf0f7;
aud[889]=16'he22f;
aud[890]=16'hd3ea;
aud[891]=16'hc666;
aud[892]=16'hb9df;
aud[893]=16'hae8b;
aud[894]=16'ha49b;
aud[895]=16'h9c3c;
aud[896]=16'h9592;
aud[897]=16'h90ba;
aud[898]=16'h8dc9;
aud[899]=16'h8ccd;
aud[900]=16'h8dc9;
aud[901]=16'h90ba;
aud[902]=16'h9592;
aud[903]=16'h9c3c;
aud[904]=16'ha49b;
aud[905]=16'hae8b;
aud[906]=16'hb9df;
aud[907]=16'hc666;
aud[908]=16'hd3ea;
aud[909]=16'he22f;
aud[910]=16'hf0f7;
aud[911]=16'h0;
aud[912]=16'hf09;
aud[913]=16'h1dd1;
aud[914]=16'h2c16;
aud[915]=16'h399a;
aud[916]=16'h4621;
aud[917]=16'h5175;
aud[918]=16'h5b65;
aud[919]=16'h63c4;
aud[920]=16'h6a6e;
aud[921]=16'h6f46;
aud[922]=16'h7237;
aud[923]=16'h7333;
aud[924]=16'h7237;
aud[925]=16'h6f46;
aud[926]=16'h6a6e;
aud[927]=16'h63c4;
aud[928]=16'h5b65;
aud[929]=16'h5175;
aud[930]=16'h4621;
aud[931]=16'h399a;
aud[932]=16'h2c16;
aud[933]=16'h1dd1;
aud[934]=16'hf09;
aud[935]=16'h0;
aud[936]=16'hf0f7;
aud[937]=16'he22f;
aud[938]=16'hd3ea;
aud[939]=16'hc666;
aud[940]=16'hb9df;
aud[941]=16'hae8b;
aud[942]=16'ha49b;
aud[943]=16'h9c3c;
aud[944]=16'h9592;
aud[945]=16'h90ba;
aud[946]=16'h8dc9;
aud[947]=16'h8ccd;
aud[948]=16'h8dc9;
aud[949]=16'h90ba;
aud[950]=16'h9592;
aud[951]=16'h9c3c;
aud[952]=16'ha49b;
aud[953]=16'hae8b;
aud[954]=16'hb9df;
aud[955]=16'hc666;
aud[956]=16'hd3ea;
aud[957]=16'he22f;
aud[958]=16'hf0f7;
aud[959]=16'h0;
aud[960]=16'hf09;
aud[961]=16'h1dd1;
aud[962]=16'h2c16;
aud[963]=16'h399a;
aud[964]=16'h4621;
aud[965]=16'h5175;
aud[966]=16'h5b65;
aud[967]=16'h63c4;
aud[968]=16'h6a6e;
aud[969]=16'h6f46;
aud[970]=16'h7237;
aud[971]=16'h7333;
aud[972]=16'h7237;
aud[973]=16'h6f46;
aud[974]=16'h6a6e;
aud[975]=16'h63c4;
aud[976]=16'h5b65;
aud[977]=16'h5175;
aud[978]=16'h4621;
aud[979]=16'h399a;
aud[980]=16'h2c16;
aud[981]=16'h1dd1;
aud[982]=16'hf09;
aud[983]=16'h0;
aud[984]=16'hf0f7;
aud[985]=16'he22f;
aud[986]=16'hd3ea;
aud[987]=16'hc666;
aud[988]=16'hb9df;
aud[989]=16'hae8b;
aud[990]=16'ha49b;
aud[991]=16'h9c3c;
aud[992]=16'h9592;
aud[993]=16'h90ba;
aud[994]=16'h8dc9;
aud[995]=16'h8ccd;
aud[996]=16'h8dc9;
aud[997]=16'h90ba;
aud[998]=16'h9592;
aud[999]=16'h9c3c;
aud[1000]=16'ha49b;
aud[1001]=16'hae8b;
aud[1002]=16'hb9df;
aud[1003]=16'hc666;
aud[1004]=16'hd3ea;
aud[1005]=16'he22f;
aud[1006]=16'hf0f7;
aud[1007]=16'h0;
aud[1008]=16'hf09;
aud[1009]=16'h1dd1;
aud[1010]=16'h2c16;
aud[1011]=16'h399a;
aud[1012]=16'h4621;
aud[1013]=16'h5175;
aud[1014]=16'h5b65;
aud[1015]=16'h63c4;
aud[1016]=16'h6a6e;
aud[1017]=16'h6f46;
aud[1018]=16'h7237;
aud[1019]=16'h7333;
aud[1020]=16'h7237;
aud[1021]=16'h6f46;
aud[1022]=16'h6a6e;
aud[1023]=16'h63c4;
aud[1024]=16'h5b65;
aud[1025]=16'h5175;
aud[1026]=16'h4621;
aud[1027]=16'h399a;
aud[1028]=16'h2c16;
aud[1029]=16'h1dd1;
aud[1030]=16'hf09;
aud[1031]=16'h0;
aud[1032]=16'hf0f7;
aud[1033]=16'he22f;
aud[1034]=16'hd3ea;
aud[1035]=16'hc666;
aud[1036]=16'hb9df;
aud[1037]=16'hae8b;
aud[1038]=16'ha49b;
aud[1039]=16'h9c3c;
aud[1040]=16'h9592;
aud[1041]=16'h90ba;
aud[1042]=16'h8dc9;
aud[1043]=16'h8ccd;
aud[1044]=16'h8dc9;
aud[1045]=16'h90ba;
aud[1046]=16'h9592;
aud[1047]=16'h9c3c;
aud[1048]=16'ha49b;
aud[1049]=16'hae8b;
aud[1050]=16'hb9df;
aud[1051]=16'hc666;
aud[1052]=16'hd3ea;
aud[1053]=16'he22f;
aud[1054]=16'hf0f7;
aud[1055]=16'h0;
aud[1056]=16'hf09;
aud[1057]=16'h1dd1;
aud[1058]=16'h2c16;
aud[1059]=16'h399a;
aud[1060]=16'h4621;
aud[1061]=16'h5175;
aud[1062]=16'h5b65;
aud[1063]=16'h63c4;
aud[1064]=16'h6a6e;
aud[1065]=16'h6f46;
aud[1066]=16'h7237;
aud[1067]=16'h7333;
aud[1068]=16'h7237;
aud[1069]=16'h6f46;
aud[1070]=16'h6a6e;
aud[1071]=16'h63c4;
aud[1072]=16'h5b65;
aud[1073]=16'h5175;
aud[1074]=16'h4621;
aud[1075]=16'h399a;
aud[1076]=16'h2c16;
aud[1077]=16'h1dd1;
aud[1078]=16'hf09;
aud[1079]=16'h0;
aud[1080]=16'hf0f7;
aud[1081]=16'he22f;
aud[1082]=16'hd3ea;
aud[1083]=16'hc666;
aud[1084]=16'hb9df;
aud[1085]=16'hae8b;
aud[1086]=16'ha49b;
aud[1087]=16'h9c3c;
aud[1088]=16'h9592;
aud[1089]=16'h90ba;
aud[1090]=16'h8dc9;
aud[1091]=16'h8ccd;
aud[1092]=16'h8dc9;
aud[1093]=16'h90ba;
aud[1094]=16'h9592;
aud[1095]=16'h9c3c;
aud[1096]=16'ha49b;
aud[1097]=16'hae8b;
aud[1098]=16'hb9df;
aud[1099]=16'hc666;
aud[1100]=16'hd3ea;
aud[1101]=16'he22f;
aud[1102]=16'hf0f7;
aud[1103]=16'h0;
aud[1104]=16'hf09;
aud[1105]=16'h1dd1;
aud[1106]=16'h2c16;
aud[1107]=16'h399a;
aud[1108]=16'h4621;
aud[1109]=16'h5175;
aud[1110]=16'h5b65;
aud[1111]=16'h63c4;
aud[1112]=16'h6a6e;
aud[1113]=16'h6f46;
aud[1114]=16'h7237;
aud[1115]=16'h7333;
aud[1116]=16'h7237;
aud[1117]=16'h6f46;
aud[1118]=16'h6a6e;
aud[1119]=16'h63c4;
aud[1120]=16'h5b65;
aud[1121]=16'h5175;
aud[1122]=16'h4621;
aud[1123]=16'h399a;
aud[1124]=16'h2c16;
aud[1125]=16'h1dd1;
aud[1126]=16'hf09;
aud[1127]=16'h0;
aud[1128]=16'hf0f7;
aud[1129]=16'he22f;
aud[1130]=16'hd3ea;
aud[1131]=16'hc666;
aud[1132]=16'hb9df;
aud[1133]=16'hae8b;
aud[1134]=16'ha49b;
aud[1135]=16'h9c3c;
aud[1136]=16'h9592;
aud[1137]=16'h90ba;
aud[1138]=16'h8dc9;
aud[1139]=16'h8ccd;
aud[1140]=16'h8dc9;
aud[1141]=16'h90ba;
aud[1142]=16'h9592;
aud[1143]=16'h9c3c;
aud[1144]=16'ha49b;
aud[1145]=16'hae8b;
aud[1146]=16'hb9df;
aud[1147]=16'hc666;
aud[1148]=16'hd3ea;
aud[1149]=16'he22f;
aud[1150]=16'hf0f7;
aud[1151]=16'h0;
aud[1152]=16'hf09;
aud[1153]=16'h1dd1;
aud[1154]=16'h2c16;
aud[1155]=16'h399a;
aud[1156]=16'h4621;
aud[1157]=16'h5175;
aud[1158]=16'h5b65;
aud[1159]=16'h63c4;
aud[1160]=16'h6a6e;
aud[1161]=16'h6f46;
aud[1162]=16'h7237;
aud[1163]=16'h7333;
aud[1164]=16'h7237;
aud[1165]=16'h6f46;
aud[1166]=16'h6a6e;
aud[1167]=16'h63c4;
aud[1168]=16'h5b65;
aud[1169]=16'h5175;
aud[1170]=16'h4621;
aud[1171]=16'h399a;
aud[1172]=16'h2c16;
aud[1173]=16'h1dd1;
aud[1174]=16'hf09;
aud[1175]=16'h0;
aud[1176]=16'hf0f7;
aud[1177]=16'he22f;
aud[1178]=16'hd3ea;
aud[1179]=16'hc666;
aud[1180]=16'hb9df;
aud[1181]=16'hae8b;
aud[1182]=16'ha49b;
aud[1183]=16'h9c3c;
aud[1184]=16'h9592;
aud[1185]=16'h90ba;
aud[1186]=16'h8dc9;
aud[1187]=16'h8ccd;
aud[1188]=16'h8dc9;
aud[1189]=16'h90ba;
aud[1190]=16'h9592;
aud[1191]=16'h9c3c;
aud[1192]=16'ha49b;
aud[1193]=16'hae8b;
aud[1194]=16'hb9df;
aud[1195]=16'hc666;
aud[1196]=16'hd3ea;
aud[1197]=16'he22f;
aud[1198]=16'hf0f7;
aud[1199]=16'h0;
aud[1200]=16'hf09;
aud[1201]=16'h1dd1;
aud[1202]=16'h2c16;
aud[1203]=16'h399a;
aud[1204]=16'h4621;
aud[1205]=16'h5175;
aud[1206]=16'h5b65;
aud[1207]=16'h63c4;
aud[1208]=16'h6a6e;
aud[1209]=16'h6f46;
aud[1210]=16'h7237;
aud[1211]=16'h7333;
aud[1212]=16'h7237;
aud[1213]=16'h6f46;
aud[1214]=16'h6a6e;
aud[1215]=16'h63c4;
aud[1216]=16'h5b65;
aud[1217]=16'h5175;
aud[1218]=16'h4621;
aud[1219]=16'h399a;
aud[1220]=16'h2c16;
aud[1221]=16'h1dd1;
aud[1222]=16'hf09;
aud[1223]=16'h0;
aud[1224]=16'hf0f7;
aud[1225]=16'he22f;
aud[1226]=16'hd3ea;
aud[1227]=16'hc666;
aud[1228]=16'hb9df;
aud[1229]=16'hae8b;
aud[1230]=16'ha49b;
aud[1231]=16'h9c3c;
aud[1232]=16'h9592;
aud[1233]=16'h90ba;
aud[1234]=16'h8dc9;
aud[1235]=16'h8ccd;
aud[1236]=16'h8dc9;
aud[1237]=16'h90ba;
aud[1238]=16'h9592;
aud[1239]=16'h9c3c;
aud[1240]=16'ha49b;
aud[1241]=16'hae8b;
aud[1242]=16'hb9df;
aud[1243]=16'hc666;
aud[1244]=16'hd3ea;
aud[1245]=16'he22f;
aud[1246]=16'hf0f7;
aud[1247]=16'h0;
aud[1248]=16'hf09;
aud[1249]=16'h1dd1;
aud[1250]=16'h2c16;
aud[1251]=16'h399a;
aud[1252]=16'h4621;
aud[1253]=16'h5175;
aud[1254]=16'h5b65;
aud[1255]=16'h63c4;
aud[1256]=16'h6a6e;
aud[1257]=16'h6f46;
aud[1258]=16'h7237;
aud[1259]=16'h7333;
aud[1260]=16'h7237;
aud[1261]=16'h6f46;
aud[1262]=16'h6a6e;
aud[1263]=16'h63c4;
aud[1264]=16'h5b65;
aud[1265]=16'h5175;
aud[1266]=16'h4621;
aud[1267]=16'h399a;
aud[1268]=16'h2c16;
aud[1269]=16'h1dd1;
aud[1270]=16'hf09;
aud[1271]=16'h0;
aud[1272]=16'hf0f7;
aud[1273]=16'he22f;
aud[1274]=16'hd3ea;
aud[1275]=16'hc666;
aud[1276]=16'hb9df;
aud[1277]=16'hae8b;
aud[1278]=16'ha49b;
aud[1279]=16'h9c3c;
aud[1280]=16'h9592;
aud[1281]=16'h90ba;
aud[1282]=16'h8dc9;
aud[1283]=16'h8ccd;
aud[1284]=16'h8dc9;
aud[1285]=16'h90ba;
aud[1286]=16'h9592;
aud[1287]=16'h9c3c;
aud[1288]=16'ha49b;
aud[1289]=16'hae8b;
aud[1290]=16'hb9df;
aud[1291]=16'hc666;
aud[1292]=16'hd3ea;
aud[1293]=16'he22f;
aud[1294]=16'hf0f7;
aud[1295]=16'h0;
aud[1296]=16'hf09;
aud[1297]=16'h1dd1;
aud[1298]=16'h2c16;
aud[1299]=16'h399a;
aud[1300]=16'h4621;
aud[1301]=16'h5175;
aud[1302]=16'h5b65;
aud[1303]=16'h63c4;
aud[1304]=16'h6a6e;
aud[1305]=16'h6f46;
aud[1306]=16'h7237;
aud[1307]=16'h7333;
aud[1308]=16'h7237;
aud[1309]=16'h6f46;
aud[1310]=16'h6a6e;
aud[1311]=16'h63c4;
aud[1312]=16'h5b65;
aud[1313]=16'h5175;
aud[1314]=16'h4621;
aud[1315]=16'h399a;
aud[1316]=16'h2c16;
aud[1317]=16'h1dd1;
aud[1318]=16'hf09;
aud[1319]=16'h0;
aud[1320]=16'hf0f7;
aud[1321]=16'he22f;
aud[1322]=16'hd3ea;
aud[1323]=16'hc666;
aud[1324]=16'hb9df;
aud[1325]=16'hae8b;
aud[1326]=16'ha49b;
aud[1327]=16'h9c3c;
aud[1328]=16'h9592;
aud[1329]=16'h90ba;
aud[1330]=16'h8dc9;
aud[1331]=16'h8ccd;
aud[1332]=16'h8dc9;
aud[1333]=16'h90ba;
aud[1334]=16'h9592;
aud[1335]=16'h9c3c;
aud[1336]=16'ha49b;
aud[1337]=16'hae8b;
aud[1338]=16'hb9df;
aud[1339]=16'hc666;
aud[1340]=16'hd3ea;
aud[1341]=16'he22f;
aud[1342]=16'hf0f7;
aud[1343]=16'h0;
aud[1344]=16'hf09;
aud[1345]=16'h1dd1;
aud[1346]=16'h2c16;
aud[1347]=16'h399a;
aud[1348]=16'h4621;
aud[1349]=16'h5175;
aud[1350]=16'h5b65;
aud[1351]=16'h63c4;
aud[1352]=16'h6a6e;
aud[1353]=16'h6f46;
aud[1354]=16'h7237;
aud[1355]=16'h7333;
aud[1356]=16'h7237;
aud[1357]=16'h6f46;
aud[1358]=16'h6a6e;
aud[1359]=16'h63c4;
aud[1360]=16'h5b65;
aud[1361]=16'h5175;
aud[1362]=16'h4621;
aud[1363]=16'h399a;
aud[1364]=16'h2c16;
aud[1365]=16'h1dd1;
aud[1366]=16'hf09;
aud[1367]=16'h0;
aud[1368]=16'hf0f7;
aud[1369]=16'he22f;
aud[1370]=16'hd3ea;
aud[1371]=16'hc666;
aud[1372]=16'hb9df;
aud[1373]=16'hae8b;
aud[1374]=16'ha49b;
aud[1375]=16'h9c3c;
aud[1376]=16'h9592;
aud[1377]=16'h90ba;
aud[1378]=16'h8dc9;
aud[1379]=16'h8ccd;
aud[1380]=16'h8dc9;
aud[1381]=16'h90ba;
aud[1382]=16'h9592;
aud[1383]=16'h9c3c;
aud[1384]=16'ha49b;
aud[1385]=16'hae8b;
aud[1386]=16'hb9df;
aud[1387]=16'hc666;
aud[1388]=16'hd3ea;
aud[1389]=16'he22f;
aud[1390]=16'hf0f7;
aud[1391]=16'h0;
aud[1392]=16'hf09;
aud[1393]=16'h1dd1;
aud[1394]=16'h2c16;
aud[1395]=16'h399a;
aud[1396]=16'h4621;
aud[1397]=16'h5175;
aud[1398]=16'h5b65;
aud[1399]=16'h63c4;
aud[1400]=16'h6a6e;
aud[1401]=16'h6f46;
aud[1402]=16'h7237;
aud[1403]=16'h7333;
aud[1404]=16'h7237;
aud[1405]=16'h6f46;
aud[1406]=16'h6a6e;
aud[1407]=16'h63c4;
aud[1408]=16'h5b65;
aud[1409]=16'h5175;
aud[1410]=16'h4621;
aud[1411]=16'h399a;
aud[1412]=16'h2c16;
aud[1413]=16'h1dd1;
aud[1414]=16'hf09;
aud[1415]=16'h0;
aud[1416]=16'hf0f7;
aud[1417]=16'he22f;
aud[1418]=16'hd3ea;
aud[1419]=16'hc666;
aud[1420]=16'hb9df;
aud[1421]=16'hae8b;
aud[1422]=16'ha49b;
aud[1423]=16'h9c3c;
aud[1424]=16'h9592;
aud[1425]=16'h90ba;
aud[1426]=16'h8dc9;
aud[1427]=16'h8ccd;
aud[1428]=16'h8dc9;
aud[1429]=16'h90ba;
aud[1430]=16'h9592;
aud[1431]=16'h9c3c;
aud[1432]=16'ha49b;
aud[1433]=16'hae8b;
aud[1434]=16'hb9df;
aud[1435]=16'hc666;
aud[1436]=16'hd3ea;
aud[1437]=16'he22f;
aud[1438]=16'hf0f7;
aud[1439]=16'h0;
aud[1440]=16'hf09;
aud[1441]=16'h1dd1;
aud[1442]=16'h2c16;
aud[1443]=16'h399a;
aud[1444]=16'h4621;
aud[1445]=16'h5175;
aud[1446]=16'h5b65;
aud[1447]=16'h63c4;
aud[1448]=16'h6a6e;
aud[1449]=16'h6f46;
aud[1450]=16'h7237;
aud[1451]=16'h7333;
aud[1452]=16'h7237;
aud[1453]=16'h6f46;
aud[1454]=16'h6a6e;
aud[1455]=16'h63c4;
aud[1456]=16'h5b65;
aud[1457]=16'h5175;
aud[1458]=16'h4621;
aud[1459]=16'h399a;
aud[1460]=16'h2c16;
aud[1461]=16'h1dd1;
aud[1462]=16'hf09;
aud[1463]=16'h0;
aud[1464]=16'hf0f7;
aud[1465]=16'he22f;
aud[1466]=16'hd3ea;
aud[1467]=16'hc666;
aud[1468]=16'hb9df;
aud[1469]=16'hae8b;
aud[1470]=16'ha49b;
aud[1471]=16'h9c3c;
aud[1472]=16'h9592;
aud[1473]=16'h90ba;
aud[1474]=16'h8dc9;
aud[1475]=16'h8ccd;
aud[1476]=16'h8dc9;
aud[1477]=16'h90ba;
aud[1478]=16'h9592;
aud[1479]=16'h9c3c;
aud[1480]=16'ha49b;
aud[1481]=16'hae8b;
aud[1482]=16'hb9df;
aud[1483]=16'hc666;
aud[1484]=16'hd3ea;
aud[1485]=16'he22f;
aud[1486]=16'hf0f7;
aud[1487]=16'h0;
aud[1488]=16'hf09;
aud[1489]=16'h1dd1;
aud[1490]=16'h2c16;
aud[1491]=16'h399a;
aud[1492]=16'h4621;
aud[1493]=16'h5175;
aud[1494]=16'h5b65;
aud[1495]=16'h63c4;
aud[1496]=16'h6a6e;
aud[1497]=16'h6f46;
aud[1498]=16'h7237;
aud[1499]=16'h7333;
aud[1500]=16'h7237;
aud[1501]=16'h6f46;
aud[1502]=16'h6a6e;
aud[1503]=16'h63c4;
aud[1504]=16'h5b65;
aud[1505]=16'h5175;
aud[1506]=16'h4621;
aud[1507]=16'h399a;
aud[1508]=16'h2c16;
aud[1509]=16'h1dd1;
aud[1510]=16'hf09;
aud[1511]=16'h0;
aud[1512]=16'hf0f7;
aud[1513]=16'he22f;
aud[1514]=16'hd3ea;
aud[1515]=16'hc666;
aud[1516]=16'hb9df;
aud[1517]=16'hae8b;
aud[1518]=16'ha49b;
aud[1519]=16'h9c3c;
aud[1520]=16'h9592;
aud[1521]=16'h90ba;
aud[1522]=16'h8dc9;
aud[1523]=16'h8ccd;
aud[1524]=16'h8dc9;
aud[1525]=16'h90ba;
aud[1526]=16'h9592;
aud[1527]=16'h9c3c;
aud[1528]=16'ha49b;
aud[1529]=16'hae8b;
aud[1530]=16'hb9df;
aud[1531]=16'hc666;
aud[1532]=16'hd3ea;
aud[1533]=16'he22f;
aud[1534]=16'hf0f7;
aud[1535]=16'h0;
aud[1536]=16'hf09;
aud[1537]=16'h1dd1;
aud[1538]=16'h2c16;
aud[1539]=16'h399a;
aud[1540]=16'h4621;
aud[1541]=16'h5175;
aud[1542]=16'h5b65;
aud[1543]=16'h63c4;
aud[1544]=16'h6a6e;
aud[1545]=16'h6f46;
aud[1546]=16'h7237;
aud[1547]=16'h7333;
aud[1548]=16'h7237;
aud[1549]=16'h6f46;
aud[1550]=16'h6a6e;
aud[1551]=16'h63c4;
aud[1552]=16'h5b65;
aud[1553]=16'h5175;
aud[1554]=16'h4621;
aud[1555]=16'h399a;
aud[1556]=16'h2c16;
aud[1557]=16'h1dd1;
aud[1558]=16'hf09;
aud[1559]=16'h0;
aud[1560]=16'hf0f7;
aud[1561]=16'he22f;
aud[1562]=16'hd3ea;
aud[1563]=16'hc666;
aud[1564]=16'hb9df;
aud[1565]=16'hae8b;
aud[1566]=16'ha49b;
aud[1567]=16'h9c3c;
aud[1568]=16'h9592;
aud[1569]=16'h90ba;
aud[1570]=16'h8dc9;
aud[1571]=16'h8ccd;
aud[1572]=16'h8dc9;
aud[1573]=16'h90ba;
aud[1574]=16'h9592;
aud[1575]=16'h9c3c;
aud[1576]=16'ha49b;
aud[1577]=16'hae8b;
aud[1578]=16'hb9df;
aud[1579]=16'hc666;
aud[1580]=16'hd3ea;
aud[1581]=16'he22f;
aud[1582]=16'hf0f7;
aud[1583]=16'h0;
aud[1584]=16'hf09;
aud[1585]=16'h1dd1;
aud[1586]=16'h2c16;
aud[1587]=16'h399a;
aud[1588]=16'h4621;
aud[1589]=16'h5175;
aud[1590]=16'h5b65;
aud[1591]=16'h63c4;
aud[1592]=16'h6a6e;
aud[1593]=16'h6f46;
aud[1594]=16'h7237;
aud[1595]=16'h7333;
aud[1596]=16'h7237;
aud[1597]=16'h6f46;
aud[1598]=16'h6a6e;
aud[1599]=16'h63c4;
aud[1600]=16'h5b65;
aud[1601]=16'h5175;
aud[1602]=16'h4621;
aud[1603]=16'h399a;
aud[1604]=16'h2c16;
aud[1605]=16'h1dd1;
aud[1606]=16'hf09;
aud[1607]=16'h0;
aud[1608]=16'hf0f7;
aud[1609]=16'he22f;
aud[1610]=16'hd3ea;
aud[1611]=16'hc666;
aud[1612]=16'hb9df;
aud[1613]=16'hae8b;
aud[1614]=16'ha49b;
aud[1615]=16'h9c3c;
aud[1616]=16'h9592;
aud[1617]=16'h90ba;
aud[1618]=16'h8dc9;
aud[1619]=16'h8ccd;
aud[1620]=16'h8dc9;
aud[1621]=16'h90ba;
aud[1622]=16'h9592;
aud[1623]=16'h9c3c;
aud[1624]=16'ha49b;
aud[1625]=16'hae8b;
aud[1626]=16'hb9df;
aud[1627]=16'hc666;
aud[1628]=16'hd3ea;
aud[1629]=16'he22f;
aud[1630]=16'hf0f7;
aud[1631]=16'h0;
aud[1632]=16'hf09;
aud[1633]=16'h1dd1;
aud[1634]=16'h2c16;
aud[1635]=16'h399a;
aud[1636]=16'h4621;
aud[1637]=16'h5175;
aud[1638]=16'h5b65;
aud[1639]=16'h63c4;
aud[1640]=16'h6a6e;
aud[1641]=16'h6f46;
aud[1642]=16'h7237;
aud[1643]=16'h7333;
aud[1644]=16'h7237;
aud[1645]=16'h6f46;
aud[1646]=16'h6a6e;
aud[1647]=16'h63c4;
aud[1648]=16'h5b65;
aud[1649]=16'h5175;
aud[1650]=16'h4621;
aud[1651]=16'h399a;
aud[1652]=16'h2c16;
aud[1653]=16'h1dd1;
aud[1654]=16'hf09;
aud[1655]=16'h0;
aud[1656]=16'hf0f7;
aud[1657]=16'he22f;
aud[1658]=16'hd3ea;
aud[1659]=16'hc666;
aud[1660]=16'hb9df;
aud[1661]=16'hae8b;
aud[1662]=16'ha49b;
aud[1663]=16'h9c3c;
aud[1664]=16'h9592;
aud[1665]=16'h90ba;
aud[1666]=16'h8dc9;
aud[1667]=16'h8ccd;
aud[1668]=16'h8dc9;
aud[1669]=16'h90ba;
aud[1670]=16'h9592;
aud[1671]=16'h9c3c;
aud[1672]=16'ha49b;
aud[1673]=16'hae8b;
aud[1674]=16'hb9df;
aud[1675]=16'hc666;
aud[1676]=16'hd3ea;
aud[1677]=16'he22f;
aud[1678]=16'hf0f7;
aud[1679]=16'h0;
aud[1680]=16'hf09;
aud[1681]=16'h1dd1;
aud[1682]=16'h2c16;
aud[1683]=16'h399a;
aud[1684]=16'h4621;
aud[1685]=16'h5175;
aud[1686]=16'h5b65;
aud[1687]=16'h63c4;
aud[1688]=16'h6a6e;
aud[1689]=16'h6f46;
aud[1690]=16'h7237;
aud[1691]=16'h7333;
aud[1692]=16'h7237;
aud[1693]=16'h6f46;
aud[1694]=16'h6a6e;
aud[1695]=16'h63c4;
aud[1696]=16'h5b65;
aud[1697]=16'h5175;
aud[1698]=16'h4621;
aud[1699]=16'h399a;
aud[1700]=16'h2c16;
aud[1701]=16'h1dd1;
aud[1702]=16'hf09;
aud[1703]=16'h0;
aud[1704]=16'hf0f7;
aud[1705]=16'he22f;
aud[1706]=16'hd3ea;
aud[1707]=16'hc666;
aud[1708]=16'hb9df;
aud[1709]=16'hae8b;
aud[1710]=16'ha49b;
aud[1711]=16'h9c3c;
aud[1712]=16'h9592;
aud[1713]=16'h90ba;
aud[1714]=16'h8dc9;
aud[1715]=16'h8ccd;
aud[1716]=16'h8dc9;
aud[1717]=16'h90ba;
aud[1718]=16'h9592;
aud[1719]=16'h9c3c;
aud[1720]=16'ha49b;
aud[1721]=16'hae8b;
aud[1722]=16'hb9df;
aud[1723]=16'hc666;
aud[1724]=16'hd3ea;
aud[1725]=16'he22f;
aud[1726]=16'hf0f7;
aud[1727]=16'h0;
aud[1728]=16'hf09;
aud[1729]=16'h1dd1;
aud[1730]=16'h2c16;
aud[1731]=16'h399a;
aud[1732]=16'h4621;
aud[1733]=16'h5175;
aud[1734]=16'h5b65;
aud[1735]=16'h63c4;
aud[1736]=16'h6a6e;
aud[1737]=16'h6f46;
aud[1738]=16'h7237;
aud[1739]=16'h7333;
aud[1740]=16'h7237;
aud[1741]=16'h6f46;
aud[1742]=16'h6a6e;
aud[1743]=16'h63c4;
aud[1744]=16'h5b65;
aud[1745]=16'h5175;
aud[1746]=16'h4621;
aud[1747]=16'h399a;
aud[1748]=16'h2c16;
aud[1749]=16'h1dd1;
aud[1750]=16'hf09;
aud[1751]=16'h0;
aud[1752]=16'hf0f7;
aud[1753]=16'he22f;
aud[1754]=16'hd3ea;
aud[1755]=16'hc666;
aud[1756]=16'hb9df;
aud[1757]=16'hae8b;
aud[1758]=16'ha49b;
aud[1759]=16'h9c3c;
aud[1760]=16'h9592;
aud[1761]=16'h90ba;
aud[1762]=16'h8dc9;
aud[1763]=16'h8ccd;
aud[1764]=16'h8dc9;
aud[1765]=16'h90ba;
aud[1766]=16'h9592;
aud[1767]=16'h9c3c;
aud[1768]=16'ha49b;
aud[1769]=16'hae8b;
aud[1770]=16'hb9df;
aud[1771]=16'hc666;
aud[1772]=16'hd3ea;
aud[1773]=16'he22f;
aud[1774]=16'hf0f7;
aud[1775]=16'h0;
aud[1776]=16'hf09;
aud[1777]=16'h1dd1;
aud[1778]=16'h2c16;
aud[1779]=16'h399a;
aud[1780]=16'h4621;
aud[1781]=16'h5175;
aud[1782]=16'h5b65;
aud[1783]=16'h63c4;
aud[1784]=16'h6a6e;
aud[1785]=16'h6f46;
aud[1786]=16'h7237;
aud[1787]=16'h7333;
aud[1788]=16'h7237;
aud[1789]=16'h6f46;
aud[1790]=16'h6a6e;
aud[1791]=16'h63c4;
aud[1792]=16'h5b65;
aud[1793]=16'h5175;
aud[1794]=16'h4621;
aud[1795]=16'h399a;
aud[1796]=16'h2c16;
aud[1797]=16'h1dd1;
aud[1798]=16'hf09;
aud[1799]=16'h0;
aud[1800]=16'hf0f7;
aud[1801]=16'he22f;
aud[1802]=16'hd3ea;
aud[1803]=16'hc666;
aud[1804]=16'hb9df;
aud[1805]=16'hae8b;
aud[1806]=16'ha49b;
aud[1807]=16'h9c3c;
aud[1808]=16'h9592;
aud[1809]=16'h90ba;
aud[1810]=16'h8dc9;
aud[1811]=16'h8ccd;
aud[1812]=16'h8dc9;
aud[1813]=16'h90ba;
aud[1814]=16'h9592;
aud[1815]=16'h9c3c;
aud[1816]=16'ha49b;
aud[1817]=16'hae8b;
aud[1818]=16'hb9df;
aud[1819]=16'hc666;
aud[1820]=16'hd3ea;
aud[1821]=16'he22f;
aud[1822]=16'hf0f7;
aud[1823]=16'h0;
aud[1824]=16'hf09;
aud[1825]=16'h1dd1;
aud[1826]=16'h2c16;
aud[1827]=16'h399a;
aud[1828]=16'h4621;
aud[1829]=16'h5175;
aud[1830]=16'h5b65;
aud[1831]=16'h63c4;
aud[1832]=16'h6a6e;
aud[1833]=16'h6f46;
aud[1834]=16'h7237;
aud[1835]=16'h7333;
aud[1836]=16'h7237;
aud[1837]=16'h6f46;
aud[1838]=16'h6a6e;
aud[1839]=16'h63c4;
aud[1840]=16'h5b65;
aud[1841]=16'h5175;
aud[1842]=16'h4621;
aud[1843]=16'h399a;
aud[1844]=16'h2c16;
aud[1845]=16'h1dd1;
aud[1846]=16'hf09;
aud[1847]=16'h0;
aud[1848]=16'hf0f7;
aud[1849]=16'he22f;
aud[1850]=16'hd3ea;
aud[1851]=16'hc666;
aud[1852]=16'hb9df;
aud[1853]=16'hae8b;
aud[1854]=16'ha49b;
aud[1855]=16'h9c3c;
aud[1856]=16'h9592;
aud[1857]=16'h90ba;
aud[1858]=16'h8dc9;
aud[1859]=16'h8ccd;
aud[1860]=16'h8dc9;
aud[1861]=16'h90ba;
aud[1862]=16'h9592;
aud[1863]=16'h9c3c;
aud[1864]=16'ha49b;
aud[1865]=16'hae8b;
aud[1866]=16'hb9df;
aud[1867]=16'hc666;
aud[1868]=16'hd3ea;
aud[1869]=16'he22f;
aud[1870]=16'hf0f7;
aud[1871]=16'h0;
aud[1872]=16'hf09;
aud[1873]=16'h1dd1;
aud[1874]=16'h2c16;
aud[1875]=16'h399a;
aud[1876]=16'h4621;
aud[1877]=16'h5175;
aud[1878]=16'h5b65;
aud[1879]=16'h63c4;
aud[1880]=16'h6a6e;
aud[1881]=16'h6f46;
aud[1882]=16'h7237;
aud[1883]=16'h7333;
aud[1884]=16'h7237;
aud[1885]=16'h6f46;
aud[1886]=16'h6a6e;
aud[1887]=16'h63c4;
aud[1888]=16'h5b65;
aud[1889]=16'h5175;
aud[1890]=16'h4621;
aud[1891]=16'h399a;
aud[1892]=16'h2c16;
aud[1893]=16'h1dd1;
aud[1894]=16'hf09;
aud[1895]=16'h0;
aud[1896]=16'hf0f7;
aud[1897]=16'he22f;
aud[1898]=16'hd3ea;
aud[1899]=16'hc666;
aud[1900]=16'hb9df;
aud[1901]=16'hae8b;
aud[1902]=16'ha49b;
aud[1903]=16'h9c3c;
aud[1904]=16'h9592;
aud[1905]=16'h90ba;
aud[1906]=16'h8dc9;
aud[1907]=16'h8ccd;
aud[1908]=16'h8dc9;
aud[1909]=16'h90ba;
aud[1910]=16'h9592;
aud[1911]=16'h9c3c;
aud[1912]=16'ha49b;
aud[1913]=16'hae8b;
aud[1914]=16'hb9df;
aud[1915]=16'hc666;
aud[1916]=16'hd3ea;
aud[1917]=16'he22f;
aud[1918]=16'hf0f7;
aud[1919]=16'h0;
aud[1920]=16'hf09;
aud[1921]=16'h1dd1;
aud[1922]=16'h2c16;
aud[1923]=16'h399a;
aud[1924]=16'h4621;
aud[1925]=16'h5175;
aud[1926]=16'h5b65;
aud[1927]=16'h63c4;
aud[1928]=16'h6a6e;
aud[1929]=16'h6f46;
aud[1930]=16'h7237;
aud[1931]=16'h7333;
aud[1932]=16'h7237;
aud[1933]=16'h6f46;
aud[1934]=16'h6a6e;
aud[1935]=16'h63c4;
aud[1936]=16'h5b65;
aud[1937]=16'h5175;
aud[1938]=16'h4621;
aud[1939]=16'h399a;
aud[1940]=16'h2c16;
aud[1941]=16'h1dd1;
aud[1942]=16'hf09;
aud[1943]=16'h0;
aud[1944]=16'hf0f7;
aud[1945]=16'he22f;
aud[1946]=16'hd3ea;
aud[1947]=16'hc666;
aud[1948]=16'hb9df;
aud[1949]=16'hae8b;
aud[1950]=16'ha49b;
aud[1951]=16'h9c3c;
aud[1952]=16'h9592;
aud[1953]=16'h90ba;
aud[1954]=16'h8dc9;
aud[1955]=16'h8ccd;
aud[1956]=16'h8dc9;
aud[1957]=16'h90ba;
aud[1958]=16'h9592;
aud[1959]=16'h9c3c;
aud[1960]=16'ha49b;
aud[1961]=16'hae8b;
aud[1962]=16'hb9df;
aud[1963]=16'hc666;
aud[1964]=16'hd3ea;
aud[1965]=16'he22f;
aud[1966]=16'hf0f7;
aud[1967]=16'h0;
aud[1968]=16'hf09;
aud[1969]=16'h1dd1;
aud[1970]=16'h2c16;
aud[1971]=16'h399a;
aud[1972]=16'h4621;
aud[1973]=16'h5175;
aud[1974]=16'h5b65;
aud[1975]=16'h63c4;
aud[1976]=16'h6a6e;
aud[1977]=16'h6f46;
aud[1978]=16'h7237;
aud[1979]=16'h7333;
aud[1980]=16'h7237;
aud[1981]=16'h6f46;
aud[1982]=16'h6a6e;
aud[1983]=16'h63c4;
aud[1984]=16'h5b65;
aud[1985]=16'h5175;
aud[1986]=16'h4621;
aud[1987]=16'h399a;
aud[1988]=16'h2c16;
aud[1989]=16'h1dd1;
aud[1990]=16'hf09;
aud[1991]=16'h0;
aud[1992]=16'hf0f7;
aud[1993]=16'he22f;
aud[1994]=16'hd3ea;
aud[1995]=16'hc666;
aud[1996]=16'hb9df;
aud[1997]=16'hae8b;
aud[1998]=16'ha49b;
aud[1999]=16'h9c3c;

end


endmodule