module testVect (
output reg signed [15:0] aud [0:1999]
);

initial begin
aud[0]=16'h2f50;
aud[1]=16'h4e62;
aud[2]=16'h539f;
aud[3]=16'h4000;
aud[4]=16'h1e9b;
aud[5]=16'h0;
aud[6]=16'hf352;
aud[7]=16'h0;
aud[8]=16'h22a3;
aud[9]=16'h4e62;
aud[10]=16'h723a;
aud[11]=16'h7fff;
aud[12]=16'h723a;
aud[13]=16'h4e62;
aud[14]=16'h22a3;
aud[15]=16'h0;
aud[16]=16'hf352;
aud[17]=16'h0;
aud[18]=16'h1e9b;
aud[19]=16'h4000;
aud[20]=16'h539f;
aud[21]=16'h4e62;
aud[22]=16'h2f50;
aud[23]=16'h0;
aud[24]=16'hd0b0;
aud[25]=16'hb19e;
aud[26]=16'hac61;
aud[27]=16'hc000;
aud[28]=16'he165;
aud[29]=16'h0;
aud[30]=16'hcae;
aud[31]=16'h0;
aud[32]=16'hdd5d;
aud[33]=16'hb19e;
aud[34]=16'h8dc6;
aud[35]=16'h8000;
aud[36]=16'h8dc6;
aud[37]=16'hb19e;
aud[38]=16'hdd5d;
aud[39]=16'h0;
aud[40]=16'hcae;
aud[41]=16'h0;
aud[42]=16'he165;
aud[43]=16'hc000;
aud[44]=16'hac61;
aud[45]=16'hb19e;
aud[46]=16'hd0b0;
aud[47]=16'h0;
aud[48]=16'h2f50;
aud[49]=16'h4e62;
aud[50]=16'h539f;
aud[51]=16'h4000;
aud[52]=16'h1e9b;
aud[53]=16'h0;
aud[54]=16'hf352;
aud[55]=16'h0;
aud[56]=16'h22a3;
aud[57]=16'h4e62;
aud[58]=16'h723a;
aud[59]=16'h7fff;
aud[60]=16'h723a;
aud[61]=16'h4e62;
aud[62]=16'h22a3;
aud[63]=16'h0;
aud[64]=16'hf352;
aud[65]=16'h0;
aud[66]=16'h1e9b;
aud[67]=16'h4000;
aud[68]=16'h539f;
aud[69]=16'h4e62;
aud[70]=16'h2f50;
aud[71]=16'h0;
aud[72]=16'hd0b0;
aud[73]=16'hb19e;
aud[74]=16'hac61;
aud[75]=16'hc000;
aud[76]=16'he165;
aud[77]=16'h0;
aud[78]=16'hcae;
aud[79]=16'h0;
aud[80]=16'hdd5d;
aud[81]=16'hb19e;
aud[82]=16'h8dc6;
aud[83]=16'h8000;
aud[84]=16'h8dc6;
aud[85]=16'hb19e;
aud[86]=16'hdd5d;
aud[87]=16'h0;
aud[88]=16'hcae;
aud[89]=16'h0;
aud[90]=16'he165;
aud[91]=16'hc000;
aud[92]=16'hac61;
aud[93]=16'hb19e;
aud[94]=16'hd0b0;
aud[95]=16'h0;
aud[96]=16'h2f50;
aud[97]=16'h4e62;
aud[98]=16'h539f;
aud[99]=16'h4000;
aud[100]=16'h1e9b;
aud[101]=16'h0;
aud[102]=16'hf352;
aud[103]=16'h0;
aud[104]=16'h22a3;
aud[105]=16'h4e62;
aud[106]=16'h723a;
aud[107]=16'h7fff;
aud[108]=16'h723a;
aud[109]=16'h4e62;
aud[110]=16'h22a3;
aud[111]=16'h0;
aud[112]=16'hf352;
aud[113]=16'h0;
aud[114]=16'h1e9b;
aud[115]=16'h4000;
aud[116]=16'h539f;
aud[117]=16'h4e62;
aud[118]=16'h2f50;
aud[119]=16'h0;
aud[120]=16'hd0b0;
aud[121]=16'hb19e;
aud[122]=16'hac61;
aud[123]=16'hc000;
aud[124]=16'he165;
aud[125]=16'h0;
aud[126]=16'hcae;
aud[127]=16'h0;
aud[128]=16'hdd5d;
aud[129]=16'hb19e;
aud[130]=16'h8dc6;
aud[131]=16'h8000;
aud[132]=16'h8dc6;
aud[133]=16'hb19e;
aud[134]=16'hdd5d;
aud[135]=16'h0;
aud[136]=16'hcae;
aud[137]=16'h0;
aud[138]=16'he165;
aud[139]=16'hc000;
aud[140]=16'hac61;
aud[141]=16'hb19e;
aud[142]=16'hd0b0;
aud[143]=16'h0;
aud[144]=16'h2f50;
aud[145]=16'h4e62;
aud[146]=16'h539f;
aud[147]=16'h4000;
aud[148]=16'h1e9b;
aud[149]=16'h0;
aud[150]=16'hf352;
aud[151]=16'h0;
aud[152]=16'h22a3;
aud[153]=16'h4e62;
aud[154]=16'h723a;
aud[155]=16'h7fff;
aud[156]=16'h723a;
aud[157]=16'h4e62;
aud[158]=16'h22a3;
aud[159]=16'h0;
aud[160]=16'hf352;
aud[161]=16'h0;
aud[162]=16'h1e9b;
aud[163]=16'h4000;
aud[164]=16'h539f;
aud[165]=16'h4e62;
aud[166]=16'h2f50;
aud[167]=16'h0;
aud[168]=16'hd0b0;
aud[169]=16'hb19e;
aud[170]=16'hac61;
aud[171]=16'hc000;
aud[172]=16'he165;
aud[173]=16'h0;
aud[174]=16'hcae;
aud[175]=16'h0;
aud[176]=16'hdd5d;
aud[177]=16'hb19e;
aud[178]=16'h8dc6;
aud[179]=16'h8000;
aud[180]=16'h8dc6;
aud[181]=16'hb19e;
aud[182]=16'hdd5d;
aud[183]=16'h0;
aud[184]=16'hcae;
aud[185]=16'h0;
aud[186]=16'he165;
aud[187]=16'hc000;
aud[188]=16'hac61;
aud[189]=16'hb19e;
aud[190]=16'hd0b0;
aud[191]=16'h0;
aud[192]=16'h2f50;
aud[193]=16'h4e62;
aud[194]=16'h539f;
aud[195]=16'h4000;
aud[196]=16'h1e9b;
aud[197]=16'h0;
aud[198]=16'hf352;
aud[199]=16'h0;
aud[200]=16'h22a3;
aud[201]=16'h4e62;
aud[202]=16'h723a;
aud[203]=16'h7fff;
aud[204]=16'h723a;
aud[205]=16'h4e62;
aud[206]=16'h22a3;
aud[207]=16'h0;
aud[208]=16'hf352;
aud[209]=16'h0;
aud[210]=16'h1e9b;
aud[211]=16'h4000;
aud[212]=16'h539f;
aud[213]=16'h4e62;
aud[214]=16'h2f50;
aud[215]=16'h0;
aud[216]=16'hd0b0;
aud[217]=16'hb19e;
aud[218]=16'hac61;
aud[219]=16'hc000;
aud[220]=16'he165;
aud[221]=16'h0;
aud[222]=16'hcae;
aud[223]=16'h0;
aud[224]=16'hdd5d;
aud[225]=16'hb19e;
aud[226]=16'h8dc6;
aud[227]=16'h8000;
aud[228]=16'h8dc6;
aud[229]=16'hb19e;
aud[230]=16'hdd5d;
aud[231]=16'h0;
aud[232]=16'hcae;
aud[233]=16'h0;
aud[234]=16'he165;
aud[235]=16'hc000;
aud[236]=16'hac61;
aud[237]=16'hb19e;
aud[238]=16'hd0b0;
aud[239]=16'h0;
aud[240]=16'h2f50;
aud[241]=16'h4e62;
aud[242]=16'h539f;
aud[243]=16'h4000;
aud[244]=16'h1e9b;
aud[245]=16'h0;
aud[246]=16'hf352;
aud[247]=16'h0;
aud[248]=16'h22a3;
aud[249]=16'h4e62;
aud[250]=16'h723a;
aud[251]=16'h7fff;
aud[252]=16'h723a;
aud[253]=16'h4e62;
aud[254]=16'h22a3;
aud[255]=16'h0;
aud[256]=16'hf352;
aud[257]=16'h0;
aud[258]=16'h1e9b;
aud[259]=16'h4000;
aud[260]=16'h539f;
aud[261]=16'h4e62;
aud[262]=16'h2f50;
aud[263]=16'h0;
aud[264]=16'hd0b0;
aud[265]=16'hb19e;
aud[266]=16'hac61;
aud[267]=16'hc000;
aud[268]=16'he165;
aud[269]=16'h0;
aud[270]=16'hcae;
aud[271]=16'h0;
aud[272]=16'hdd5d;
aud[273]=16'hb19e;
aud[274]=16'h8dc6;
aud[275]=16'h8000;
aud[276]=16'h8dc6;
aud[277]=16'hb19e;
aud[278]=16'hdd5d;
aud[279]=16'h0;
aud[280]=16'hcae;
aud[281]=16'h0;
aud[282]=16'he165;
aud[283]=16'hc000;
aud[284]=16'hac61;
aud[285]=16'hb19e;
aud[286]=16'hd0b0;
aud[287]=16'h0;
aud[288]=16'h2f50;
aud[289]=16'h4e62;
aud[290]=16'h539f;
aud[291]=16'h4000;
aud[292]=16'h1e9b;
aud[293]=16'h0;
aud[294]=16'hf352;
aud[295]=16'h0;
aud[296]=16'h22a3;
aud[297]=16'h4e62;
aud[298]=16'h723a;
aud[299]=16'h7fff;
aud[300]=16'h723a;
aud[301]=16'h4e62;
aud[302]=16'h22a3;
aud[303]=16'h0;
aud[304]=16'hf352;
aud[305]=16'h0;
aud[306]=16'h1e9b;
aud[307]=16'h4000;
aud[308]=16'h539f;
aud[309]=16'h4e62;
aud[310]=16'h2f50;
aud[311]=16'h0;
aud[312]=16'hd0b0;
aud[313]=16'hb19e;
aud[314]=16'hac61;
aud[315]=16'hc000;
aud[316]=16'he165;
aud[317]=16'h0;
aud[318]=16'hcae;
aud[319]=16'h0;
aud[320]=16'hdd5d;
aud[321]=16'hb19e;
aud[322]=16'h8dc6;
aud[323]=16'h8000;
aud[324]=16'h8dc6;
aud[325]=16'hb19e;
aud[326]=16'hdd5d;
aud[327]=16'h0;
aud[328]=16'hcae;
aud[329]=16'h0;
aud[330]=16'he165;
aud[331]=16'hc000;
aud[332]=16'hac61;
aud[333]=16'hb19e;
aud[334]=16'hd0b0;
aud[335]=16'h0;
aud[336]=16'h2f50;
aud[337]=16'h4e62;
aud[338]=16'h539f;
aud[339]=16'h4000;
aud[340]=16'h1e9b;
aud[341]=16'h0;
aud[342]=16'hf352;
aud[343]=16'h0;
aud[344]=16'h22a3;
aud[345]=16'h4e62;
aud[346]=16'h723a;
aud[347]=16'h7fff;
aud[348]=16'h723a;
aud[349]=16'h4e62;
aud[350]=16'h22a3;
aud[351]=16'h0;
aud[352]=16'hf352;
aud[353]=16'h0;
aud[354]=16'h1e9b;
aud[355]=16'h4000;
aud[356]=16'h539f;
aud[357]=16'h4e62;
aud[358]=16'h2f50;
aud[359]=16'h0;
aud[360]=16'hd0b0;
aud[361]=16'hb19e;
aud[362]=16'hac61;
aud[363]=16'hc000;
aud[364]=16'he165;
aud[365]=16'h0;
aud[366]=16'hcae;
aud[367]=16'h0;
aud[368]=16'hdd5d;
aud[369]=16'hb19e;
aud[370]=16'h8dc6;
aud[371]=16'h8000;
aud[372]=16'h8dc6;
aud[373]=16'hb19e;
aud[374]=16'hdd5d;
aud[375]=16'h0;
aud[376]=16'hcae;
aud[377]=16'h0;
aud[378]=16'he165;
aud[379]=16'hc000;
aud[380]=16'hac61;
aud[381]=16'hb19e;
aud[382]=16'hd0b0;
aud[383]=16'h0;
aud[384]=16'h2f50;
aud[385]=16'h4e62;
aud[386]=16'h539f;
aud[387]=16'h4000;
aud[388]=16'h1e9b;
aud[389]=16'h0;
aud[390]=16'hf352;
aud[391]=16'h0;
aud[392]=16'h22a3;
aud[393]=16'h4e62;
aud[394]=16'h723a;
aud[395]=16'h7fff;
aud[396]=16'h723a;
aud[397]=16'h4e62;
aud[398]=16'h22a3;
aud[399]=16'h0;
aud[400]=16'hf352;
aud[401]=16'h0;
aud[402]=16'h1e9b;
aud[403]=16'h4000;
aud[404]=16'h539f;
aud[405]=16'h4e62;
aud[406]=16'h2f50;
aud[407]=16'h0;
aud[408]=16'hd0b0;
aud[409]=16'hb19e;
aud[410]=16'hac61;
aud[411]=16'hc000;
aud[412]=16'he165;
aud[413]=16'h0;
aud[414]=16'hcae;
aud[415]=16'h0;
aud[416]=16'hdd5d;
aud[417]=16'hb19e;
aud[418]=16'h8dc6;
aud[419]=16'h8000;
aud[420]=16'h8dc6;
aud[421]=16'hb19e;
aud[422]=16'hdd5d;
aud[423]=16'h0;
aud[424]=16'hcae;
aud[425]=16'h0;
aud[426]=16'he165;
aud[427]=16'hc000;
aud[428]=16'hac61;
aud[429]=16'hb19e;
aud[430]=16'hd0b0;
aud[431]=16'h0;
aud[432]=16'h2f50;
aud[433]=16'h4e62;
aud[434]=16'h539f;
aud[435]=16'h4000;
aud[436]=16'h1e9b;
aud[437]=16'h0;
aud[438]=16'hf352;
aud[439]=16'h0;
aud[440]=16'h22a3;
aud[441]=16'h4e62;
aud[442]=16'h723a;
aud[443]=16'h7fff;
aud[444]=16'h723a;
aud[445]=16'h4e62;
aud[446]=16'h22a3;
aud[447]=16'h0;
aud[448]=16'hf352;
aud[449]=16'h0;
aud[450]=16'h1e9b;
aud[451]=16'h4000;
aud[452]=16'h539f;
aud[453]=16'h4e62;
aud[454]=16'h2f50;
aud[455]=16'h0;
aud[456]=16'hd0b0;
aud[457]=16'hb19e;
aud[458]=16'hac61;
aud[459]=16'hc000;
aud[460]=16'he165;
aud[461]=16'h0;
aud[462]=16'hcae;
aud[463]=16'h0;
aud[464]=16'hdd5d;
aud[465]=16'hb19e;
aud[466]=16'h8dc6;
aud[467]=16'h8000;
aud[468]=16'h8dc6;
aud[469]=16'hb19e;
aud[470]=16'hdd5d;
aud[471]=16'h0;
aud[472]=16'hcae;
aud[473]=16'h0;
aud[474]=16'he165;
aud[475]=16'hc000;
aud[476]=16'hac61;
aud[477]=16'hb19e;
aud[478]=16'hd0b0;
aud[479]=16'h0;
aud[480]=16'h2f50;
aud[481]=16'h4e62;
aud[482]=16'h539f;
aud[483]=16'h4000;
aud[484]=16'h1e9b;
aud[485]=16'h0;
aud[486]=16'hf352;
aud[487]=16'h0;
aud[488]=16'h22a3;
aud[489]=16'h4e62;
aud[490]=16'h723a;
aud[491]=16'h7fff;
aud[492]=16'h723a;
aud[493]=16'h4e62;
aud[494]=16'h22a3;
aud[495]=16'h0;
aud[496]=16'hf352;
aud[497]=16'h0;
aud[498]=16'h1e9b;
aud[499]=16'h4000;
aud[500]=16'h539f;
aud[501]=16'h4e62;
aud[502]=16'h2f50;
aud[503]=16'h0;
aud[504]=16'hd0b0;
aud[505]=16'hb19e;
aud[506]=16'hac61;
aud[507]=16'hc000;
aud[508]=16'he165;
aud[509]=16'h0;
aud[510]=16'hcae;
aud[511]=16'h0;
aud[512]=16'hdd5d;
aud[513]=16'hb19e;
aud[514]=16'h8dc6;
aud[515]=16'h8000;
aud[516]=16'h8dc6;
aud[517]=16'hb19e;
aud[518]=16'hdd5d;
aud[519]=16'h0;
aud[520]=16'hcae;
aud[521]=16'h0;
aud[522]=16'he165;
aud[523]=16'hc000;
aud[524]=16'hac61;
aud[525]=16'hb19e;
aud[526]=16'hd0b0;
aud[527]=16'h0;
aud[528]=16'h2f50;
aud[529]=16'h4e62;
aud[530]=16'h539f;
aud[531]=16'h4000;
aud[532]=16'h1e9b;
aud[533]=16'h0;
aud[534]=16'hf352;
aud[535]=16'h0;
aud[536]=16'h22a3;
aud[537]=16'h4e62;
aud[538]=16'h723a;
aud[539]=16'h7fff;
aud[540]=16'h723a;
aud[541]=16'h4e62;
aud[542]=16'h22a3;
aud[543]=16'h0;
aud[544]=16'hf352;
aud[545]=16'h0;
aud[546]=16'h1e9b;
aud[547]=16'h4000;
aud[548]=16'h539f;
aud[549]=16'h4e62;
aud[550]=16'h2f50;
aud[551]=16'h0;
aud[552]=16'hd0b0;
aud[553]=16'hb19e;
aud[554]=16'hac61;
aud[555]=16'hc000;
aud[556]=16'he165;
aud[557]=16'h0;
aud[558]=16'hcae;
aud[559]=16'h0;
aud[560]=16'hdd5d;
aud[561]=16'hb19e;
aud[562]=16'h8dc6;
aud[563]=16'h8000;
aud[564]=16'h8dc6;
aud[565]=16'hb19e;
aud[566]=16'hdd5d;
aud[567]=16'h0;
aud[568]=16'hcae;
aud[569]=16'h0;
aud[570]=16'he165;
aud[571]=16'hc000;
aud[572]=16'hac61;
aud[573]=16'hb19e;
aud[574]=16'hd0b0;
aud[575]=16'h0;
aud[576]=16'h2f50;
aud[577]=16'h4e62;
aud[578]=16'h539f;
aud[579]=16'h4000;
aud[580]=16'h1e9b;
aud[581]=16'h0;
aud[582]=16'hf352;
aud[583]=16'h0;
aud[584]=16'h22a3;
aud[585]=16'h4e62;
aud[586]=16'h723a;
aud[587]=16'h7fff;
aud[588]=16'h723a;
aud[589]=16'h4e62;
aud[590]=16'h22a3;
aud[591]=16'h0;
aud[592]=16'hf352;
aud[593]=16'h0;
aud[594]=16'h1e9b;
aud[595]=16'h4000;
aud[596]=16'h539f;
aud[597]=16'h4e62;
aud[598]=16'h2f50;
aud[599]=16'h0;
aud[600]=16'hd0b0;
aud[601]=16'hb19e;
aud[602]=16'hac61;
aud[603]=16'hc000;
aud[604]=16'he165;
aud[605]=16'h0;
aud[606]=16'hcae;
aud[607]=16'h0;
aud[608]=16'hdd5d;
aud[609]=16'hb19e;
aud[610]=16'h8dc6;
aud[611]=16'h8000;
aud[612]=16'h8dc6;
aud[613]=16'hb19e;
aud[614]=16'hdd5d;
aud[615]=16'h0;
aud[616]=16'hcae;
aud[617]=16'h0;
aud[618]=16'he165;
aud[619]=16'hc000;
aud[620]=16'hac61;
aud[621]=16'hb19e;
aud[622]=16'hd0b0;
aud[623]=16'h0;
aud[624]=16'h2f50;
aud[625]=16'h4e62;
aud[626]=16'h539f;
aud[627]=16'h4000;
aud[628]=16'h1e9b;
aud[629]=16'h0;
aud[630]=16'hf352;
aud[631]=16'h0;
aud[632]=16'h22a3;
aud[633]=16'h4e62;
aud[634]=16'h723a;
aud[635]=16'h7fff;
aud[636]=16'h723a;
aud[637]=16'h4e62;
aud[638]=16'h22a3;
aud[639]=16'h0;
aud[640]=16'hf352;
aud[641]=16'h0;
aud[642]=16'h1e9b;
aud[643]=16'h4000;
aud[644]=16'h539f;
aud[645]=16'h4e62;
aud[646]=16'h2f50;
aud[647]=16'h0;
aud[648]=16'hd0b0;
aud[649]=16'hb19e;
aud[650]=16'hac61;
aud[651]=16'hc000;
aud[652]=16'he165;
aud[653]=16'h0;
aud[654]=16'hcae;
aud[655]=16'h0;
aud[656]=16'hdd5d;
aud[657]=16'hb19e;
aud[658]=16'h8dc6;
aud[659]=16'h8000;
aud[660]=16'h8dc6;
aud[661]=16'hb19e;
aud[662]=16'hdd5d;
aud[663]=16'h0;
aud[664]=16'hcae;
aud[665]=16'h0;
aud[666]=16'he165;
aud[667]=16'hc000;
aud[668]=16'hac61;
aud[669]=16'hb19e;
aud[670]=16'hd0b0;
aud[671]=16'h0;
aud[672]=16'h2f50;
aud[673]=16'h4e62;
aud[674]=16'h539f;
aud[675]=16'h4000;
aud[676]=16'h1e9b;
aud[677]=16'h0;
aud[678]=16'hf352;
aud[679]=16'h0;
aud[680]=16'h22a3;
aud[681]=16'h4e62;
aud[682]=16'h723a;
aud[683]=16'h7fff;
aud[684]=16'h723a;
aud[685]=16'h4e62;
aud[686]=16'h22a3;
aud[687]=16'h0;
aud[688]=16'hf352;
aud[689]=16'h0;
aud[690]=16'h1e9b;
aud[691]=16'h4000;
aud[692]=16'h539f;
aud[693]=16'h4e62;
aud[694]=16'h2f50;
aud[695]=16'h0;
aud[696]=16'hd0b0;
aud[697]=16'hb19e;
aud[698]=16'hac61;
aud[699]=16'hc000;
aud[700]=16'he165;
aud[701]=16'h0;
aud[702]=16'hcae;
aud[703]=16'h0;
aud[704]=16'hdd5d;
aud[705]=16'hb19e;
aud[706]=16'h8dc6;
aud[707]=16'h8000;
aud[708]=16'h8dc6;
aud[709]=16'hb19e;
aud[710]=16'hdd5d;
aud[711]=16'h0;
aud[712]=16'hcae;
aud[713]=16'h0;
aud[714]=16'he165;
aud[715]=16'hc000;
aud[716]=16'hac61;
aud[717]=16'hb19e;
aud[718]=16'hd0b0;
aud[719]=16'h0;
aud[720]=16'h2f50;
aud[721]=16'h4e62;
aud[722]=16'h539f;
aud[723]=16'h4000;
aud[724]=16'h1e9b;
aud[725]=16'h0;
aud[726]=16'hf352;
aud[727]=16'h0;
aud[728]=16'h22a3;
aud[729]=16'h4e62;
aud[730]=16'h723a;
aud[731]=16'h7fff;
aud[732]=16'h723a;
aud[733]=16'h4e62;
aud[734]=16'h22a3;
aud[735]=16'h0;
aud[736]=16'hf352;
aud[737]=16'h0;
aud[738]=16'h1e9b;
aud[739]=16'h4000;
aud[740]=16'h539f;
aud[741]=16'h4e62;
aud[742]=16'h2f50;
aud[743]=16'h0;
aud[744]=16'hd0b0;
aud[745]=16'hb19e;
aud[746]=16'hac61;
aud[747]=16'hc000;
aud[748]=16'he165;
aud[749]=16'h0;
aud[750]=16'hcae;
aud[751]=16'h0;
aud[752]=16'hdd5d;
aud[753]=16'hb19e;
aud[754]=16'h8dc6;
aud[755]=16'h8000;
aud[756]=16'h8dc6;
aud[757]=16'hb19e;
aud[758]=16'hdd5d;
aud[759]=16'h0;
aud[760]=16'hcae;
aud[761]=16'h0;
aud[762]=16'he165;
aud[763]=16'hc000;
aud[764]=16'hac61;
aud[765]=16'hb19e;
aud[766]=16'hd0b0;
aud[767]=16'h0;
aud[768]=16'h2f50;
aud[769]=16'h4e62;
aud[770]=16'h539f;
aud[771]=16'h4000;
aud[772]=16'h1e9b;
aud[773]=16'h0;
aud[774]=16'hf352;
aud[775]=16'h0;
aud[776]=16'h22a3;
aud[777]=16'h4e62;
aud[778]=16'h723a;
aud[779]=16'h7fff;
aud[780]=16'h723a;
aud[781]=16'h4e62;
aud[782]=16'h22a3;
aud[783]=16'h0;
aud[784]=16'hf352;
aud[785]=16'h0;
aud[786]=16'h1e9b;
aud[787]=16'h4000;
aud[788]=16'h539f;
aud[789]=16'h4e62;
aud[790]=16'h2f50;
aud[791]=16'h0;
aud[792]=16'hd0b0;
aud[793]=16'hb19e;
aud[794]=16'hac61;
aud[795]=16'hc000;
aud[796]=16'he165;
aud[797]=16'h0;
aud[798]=16'hcae;
aud[799]=16'h0;
aud[800]=16'hdd5d;
aud[801]=16'hb19e;
aud[802]=16'h8dc6;
aud[803]=16'h8000;
aud[804]=16'h8dc6;
aud[805]=16'hb19e;
aud[806]=16'hdd5d;
aud[807]=16'h0;
aud[808]=16'hcae;
aud[809]=16'h0;
aud[810]=16'he165;
aud[811]=16'hc000;
aud[812]=16'hac61;
aud[813]=16'hb19e;
aud[814]=16'hd0b0;
aud[815]=16'h0;
aud[816]=16'h2f50;
aud[817]=16'h4e62;
aud[818]=16'h539f;
aud[819]=16'h4000;
aud[820]=16'h1e9b;
aud[821]=16'h0;
aud[822]=16'hf352;
aud[823]=16'h0;
aud[824]=16'h22a3;
aud[825]=16'h4e62;
aud[826]=16'h723a;
aud[827]=16'h7fff;
aud[828]=16'h723a;
aud[829]=16'h4e62;
aud[830]=16'h22a3;
aud[831]=16'h0;
aud[832]=16'hf352;
aud[833]=16'h0;
aud[834]=16'h1e9b;
aud[835]=16'h4000;
aud[836]=16'h539f;
aud[837]=16'h4e62;
aud[838]=16'h2f50;
aud[839]=16'h0;
aud[840]=16'hd0b0;
aud[841]=16'hb19e;
aud[842]=16'hac61;
aud[843]=16'hc000;
aud[844]=16'he165;
aud[845]=16'h0;
aud[846]=16'hcae;
aud[847]=16'h0;
aud[848]=16'hdd5d;
aud[849]=16'hb19e;
aud[850]=16'h8dc6;
aud[851]=16'h8000;
aud[852]=16'h8dc6;
aud[853]=16'hb19e;
aud[854]=16'hdd5d;
aud[855]=16'h0;
aud[856]=16'hcae;
aud[857]=16'h0;
aud[858]=16'he165;
aud[859]=16'hc000;
aud[860]=16'hac61;
aud[861]=16'hb19e;
aud[862]=16'hd0b0;
aud[863]=16'h0;
aud[864]=16'h2f50;
aud[865]=16'h4e62;
aud[866]=16'h539f;
aud[867]=16'h4000;
aud[868]=16'h1e9b;
aud[869]=16'h0;
aud[870]=16'hf352;
aud[871]=16'h0;
aud[872]=16'h22a3;
aud[873]=16'h4e62;
aud[874]=16'h723a;
aud[875]=16'h7fff;
aud[876]=16'h723a;
aud[877]=16'h4e62;
aud[878]=16'h22a3;
aud[879]=16'h0;
aud[880]=16'hf352;
aud[881]=16'h0;
aud[882]=16'h1e9b;
aud[883]=16'h4000;
aud[884]=16'h539f;
aud[885]=16'h4e62;
aud[886]=16'h2f50;
aud[887]=16'h0;
aud[888]=16'hd0b0;
aud[889]=16'hb19e;
aud[890]=16'hac61;
aud[891]=16'hc000;
aud[892]=16'he165;
aud[893]=16'h0;
aud[894]=16'hcae;
aud[895]=16'h0;
aud[896]=16'hdd5d;
aud[897]=16'hb19e;
aud[898]=16'h8dc6;
aud[899]=16'h8000;
aud[900]=16'h8dc6;
aud[901]=16'hb19e;
aud[902]=16'hdd5d;
aud[903]=16'h0;
aud[904]=16'hcae;
aud[905]=16'h0;
aud[906]=16'he165;
aud[907]=16'hc000;
aud[908]=16'hac61;
aud[909]=16'hb19e;
aud[910]=16'hd0b0;
aud[911]=16'h0;
aud[912]=16'h2f50;
aud[913]=16'h4e62;
aud[914]=16'h539f;
aud[915]=16'h4000;
aud[916]=16'h1e9b;
aud[917]=16'h0;
aud[918]=16'hf352;
aud[919]=16'h0;
aud[920]=16'h22a3;
aud[921]=16'h4e62;
aud[922]=16'h723a;
aud[923]=16'h7fff;
aud[924]=16'h723a;
aud[925]=16'h4e62;
aud[926]=16'h22a3;
aud[927]=16'h0;
aud[928]=16'hf352;
aud[929]=16'h0;
aud[930]=16'h1e9b;
aud[931]=16'h4000;
aud[932]=16'h539f;
aud[933]=16'h4e62;
aud[934]=16'h2f50;
aud[935]=16'h0;
aud[936]=16'hd0b0;
aud[937]=16'hb19e;
aud[938]=16'hac61;
aud[939]=16'hc000;
aud[940]=16'he165;
aud[941]=16'h0;
aud[942]=16'hcae;
aud[943]=16'h0;
aud[944]=16'hdd5d;
aud[945]=16'hb19e;
aud[946]=16'h8dc6;
aud[947]=16'h8000;
aud[948]=16'h8dc6;
aud[949]=16'hb19e;
aud[950]=16'hdd5d;
aud[951]=16'h0;
aud[952]=16'hcae;
aud[953]=16'h0;
aud[954]=16'he165;
aud[955]=16'hc000;
aud[956]=16'hac61;
aud[957]=16'hb19e;
aud[958]=16'hd0b0;
aud[959]=16'h0;
aud[960]=16'h2f50;
aud[961]=16'h4e62;
aud[962]=16'h539f;
aud[963]=16'h4000;
aud[964]=16'h1e9b;
aud[965]=16'h0;
aud[966]=16'hf352;
aud[967]=16'h0;
aud[968]=16'h22a3;
aud[969]=16'h4e62;
aud[970]=16'h723a;
aud[971]=16'h7fff;
aud[972]=16'h723a;
aud[973]=16'h4e62;
aud[974]=16'h22a3;
aud[975]=16'h0;
aud[976]=16'hf352;
aud[977]=16'h0;
aud[978]=16'h1e9b;
aud[979]=16'h4000;
aud[980]=16'h539f;
aud[981]=16'h4e62;
aud[982]=16'h2f50;
aud[983]=16'h0;
aud[984]=16'hd0b0;
aud[985]=16'hb19e;
aud[986]=16'hac61;
aud[987]=16'hc000;
aud[988]=16'he165;
aud[989]=16'h0;
aud[990]=16'hcae;
aud[991]=16'h0;
aud[992]=16'hdd5d;
aud[993]=16'hb19e;
aud[994]=16'h8dc6;
aud[995]=16'h8000;
aud[996]=16'h8dc6;
aud[997]=16'hb19e;
aud[998]=16'hdd5d;
aud[999]=16'h0;
aud[1000]=16'hcae;
aud[1001]=16'h0;
aud[1002]=16'he165;
aud[1003]=16'hc000;
aud[1004]=16'hac61;
aud[1005]=16'hb19e;
aud[1006]=16'hd0b0;
aud[1007]=16'h0;
aud[1008]=16'h2f50;
aud[1009]=16'h4e62;
aud[1010]=16'h539f;
aud[1011]=16'h4000;
aud[1012]=16'h1e9b;
aud[1013]=16'h0;
aud[1014]=16'hf352;
aud[1015]=16'h0;
aud[1016]=16'h22a3;
aud[1017]=16'h4e62;
aud[1018]=16'h723a;
aud[1019]=16'h7fff;
aud[1020]=16'h723a;
aud[1021]=16'h4e62;
aud[1022]=16'h22a3;
aud[1023]=16'h0;
aud[1024]=16'hf352;
aud[1025]=16'h0;
aud[1026]=16'h1e9b;
aud[1027]=16'h4000;
aud[1028]=16'h539f;
aud[1029]=16'h4e62;
aud[1030]=16'h2f50;
aud[1031]=16'h0;
aud[1032]=16'hd0b0;
aud[1033]=16'hb19e;
aud[1034]=16'hac61;
aud[1035]=16'hc000;
aud[1036]=16'he165;
aud[1037]=16'h0;
aud[1038]=16'hcae;
aud[1039]=16'h0;
aud[1040]=16'hdd5d;
aud[1041]=16'hb19e;
aud[1042]=16'h8dc6;
aud[1043]=16'h8000;
aud[1044]=16'h8dc6;
aud[1045]=16'hb19e;
aud[1046]=16'hdd5d;
aud[1047]=16'h0;
aud[1048]=16'hcae;
aud[1049]=16'h0;
aud[1050]=16'he165;
aud[1051]=16'hc000;
aud[1052]=16'hac61;
aud[1053]=16'hb19e;
aud[1054]=16'hd0b0;
aud[1055]=16'h0;
aud[1056]=16'h2f50;
aud[1057]=16'h4e62;
aud[1058]=16'h539f;
aud[1059]=16'h4000;
aud[1060]=16'h1e9b;
aud[1061]=16'h0;
aud[1062]=16'hf352;
aud[1063]=16'h0;
aud[1064]=16'h22a3;
aud[1065]=16'h4e62;
aud[1066]=16'h723a;
aud[1067]=16'h7fff;
aud[1068]=16'h723a;
aud[1069]=16'h4e62;
aud[1070]=16'h22a3;
aud[1071]=16'h0;
aud[1072]=16'hf352;
aud[1073]=16'h0;
aud[1074]=16'h1e9b;
aud[1075]=16'h4000;
aud[1076]=16'h539f;
aud[1077]=16'h4e62;
aud[1078]=16'h2f50;
aud[1079]=16'h0;
aud[1080]=16'hd0b0;
aud[1081]=16'hb19e;
aud[1082]=16'hac61;
aud[1083]=16'hc000;
aud[1084]=16'he165;
aud[1085]=16'h0;
aud[1086]=16'hcae;
aud[1087]=16'h0;
aud[1088]=16'hdd5d;
aud[1089]=16'hb19e;
aud[1090]=16'h8dc6;
aud[1091]=16'h8000;
aud[1092]=16'h8dc6;
aud[1093]=16'hb19e;
aud[1094]=16'hdd5d;
aud[1095]=16'h0;
aud[1096]=16'hcae;
aud[1097]=16'h0;
aud[1098]=16'he165;
aud[1099]=16'hc000;
aud[1100]=16'hac61;
aud[1101]=16'hb19e;
aud[1102]=16'hd0b0;
aud[1103]=16'h0;
aud[1104]=16'h2f50;
aud[1105]=16'h4e62;
aud[1106]=16'h539f;
aud[1107]=16'h4000;
aud[1108]=16'h1e9b;
aud[1109]=16'h0;
aud[1110]=16'hf352;
aud[1111]=16'h0;
aud[1112]=16'h22a3;
aud[1113]=16'h4e62;
aud[1114]=16'h723a;
aud[1115]=16'h7fff;
aud[1116]=16'h723a;
aud[1117]=16'h4e62;
aud[1118]=16'h22a3;
aud[1119]=16'h0;
aud[1120]=16'hf352;
aud[1121]=16'h0;
aud[1122]=16'h1e9b;
aud[1123]=16'h4000;
aud[1124]=16'h539f;
aud[1125]=16'h4e62;
aud[1126]=16'h2f50;
aud[1127]=16'h0;
aud[1128]=16'hd0b0;
aud[1129]=16'hb19e;
aud[1130]=16'hac61;
aud[1131]=16'hc000;
aud[1132]=16'he165;
aud[1133]=16'h0;
aud[1134]=16'hcae;
aud[1135]=16'h0;
aud[1136]=16'hdd5d;
aud[1137]=16'hb19e;
aud[1138]=16'h8dc6;
aud[1139]=16'h8000;
aud[1140]=16'h8dc6;
aud[1141]=16'hb19e;
aud[1142]=16'hdd5d;
aud[1143]=16'h0;
aud[1144]=16'hcae;
aud[1145]=16'h0;
aud[1146]=16'he165;
aud[1147]=16'hc000;
aud[1148]=16'hac61;
aud[1149]=16'hb19e;
aud[1150]=16'hd0b0;
aud[1151]=16'h0;
aud[1152]=16'h2f50;
aud[1153]=16'h4e62;
aud[1154]=16'h539f;
aud[1155]=16'h4000;
aud[1156]=16'h1e9b;
aud[1157]=16'h0;
aud[1158]=16'hf352;
aud[1159]=16'h0;
aud[1160]=16'h22a3;
aud[1161]=16'h4e62;
aud[1162]=16'h723a;
aud[1163]=16'h7fff;
aud[1164]=16'h723a;
aud[1165]=16'h4e62;
aud[1166]=16'h22a3;
aud[1167]=16'h0;
aud[1168]=16'hf352;
aud[1169]=16'h0;
aud[1170]=16'h1e9b;
aud[1171]=16'h4000;
aud[1172]=16'h539f;
aud[1173]=16'h4e62;
aud[1174]=16'h2f50;
aud[1175]=16'h0;
aud[1176]=16'hd0b0;
aud[1177]=16'hb19e;
aud[1178]=16'hac61;
aud[1179]=16'hc000;
aud[1180]=16'he165;
aud[1181]=16'h0;
aud[1182]=16'hcae;
aud[1183]=16'h0;
aud[1184]=16'hdd5d;
aud[1185]=16'hb19e;
aud[1186]=16'h8dc6;
aud[1187]=16'h8000;
aud[1188]=16'h8dc6;
aud[1189]=16'hb19e;
aud[1190]=16'hdd5d;
aud[1191]=16'h0;
aud[1192]=16'hcae;
aud[1193]=16'h0;
aud[1194]=16'he165;
aud[1195]=16'hc000;
aud[1196]=16'hac61;
aud[1197]=16'hb19e;
aud[1198]=16'hd0b0;
aud[1199]=16'h0;
aud[1200]=16'h2f50;
aud[1201]=16'h4e62;
aud[1202]=16'h539f;
aud[1203]=16'h4000;
aud[1204]=16'h1e9b;
aud[1205]=16'h0;
aud[1206]=16'hf352;
aud[1207]=16'h0;
aud[1208]=16'h22a3;
aud[1209]=16'h4e62;
aud[1210]=16'h723a;
aud[1211]=16'h7fff;
aud[1212]=16'h723a;
aud[1213]=16'h4e62;
aud[1214]=16'h22a3;
aud[1215]=16'h0;
aud[1216]=16'hf352;
aud[1217]=16'h0;
aud[1218]=16'h1e9b;
aud[1219]=16'h4000;
aud[1220]=16'h539f;
aud[1221]=16'h4e62;
aud[1222]=16'h2f50;
aud[1223]=16'h0;
aud[1224]=16'hd0b0;
aud[1225]=16'hb19e;
aud[1226]=16'hac61;
aud[1227]=16'hc000;
aud[1228]=16'he165;
aud[1229]=16'h0;
aud[1230]=16'hcae;
aud[1231]=16'h0;
aud[1232]=16'hdd5d;
aud[1233]=16'hb19e;
aud[1234]=16'h8dc6;
aud[1235]=16'h8000;
aud[1236]=16'h8dc6;
aud[1237]=16'hb19e;
aud[1238]=16'hdd5d;
aud[1239]=16'h0;
aud[1240]=16'hcae;
aud[1241]=16'h0;
aud[1242]=16'he165;
aud[1243]=16'hc000;
aud[1244]=16'hac61;
aud[1245]=16'hb19e;
aud[1246]=16'hd0b0;
aud[1247]=16'h0;
aud[1248]=16'h2f50;
aud[1249]=16'h4e62;
aud[1250]=16'h539f;
aud[1251]=16'h4000;
aud[1252]=16'h1e9b;
aud[1253]=16'h0;
aud[1254]=16'hf352;
aud[1255]=16'h0;
aud[1256]=16'h22a3;
aud[1257]=16'h4e62;
aud[1258]=16'h723a;
aud[1259]=16'h7fff;
aud[1260]=16'h723a;
aud[1261]=16'h4e62;
aud[1262]=16'h22a3;
aud[1263]=16'h0;
aud[1264]=16'hf352;
aud[1265]=16'h0;
aud[1266]=16'h1e9b;
aud[1267]=16'h4000;
aud[1268]=16'h539f;
aud[1269]=16'h4e62;
aud[1270]=16'h2f50;
aud[1271]=16'h0;
aud[1272]=16'hd0b0;
aud[1273]=16'hb19e;
aud[1274]=16'hac61;
aud[1275]=16'hc000;
aud[1276]=16'he165;
aud[1277]=16'h0;
aud[1278]=16'hcae;
aud[1279]=16'h0;
aud[1280]=16'hdd5d;
aud[1281]=16'hb19e;
aud[1282]=16'h8dc6;
aud[1283]=16'h8000;
aud[1284]=16'h8dc6;
aud[1285]=16'hb19e;
aud[1286]=16'hdd5d;
aud[1287]=16'h0;
aud[1288]=16'hcae;
aud[1289]=16'h0;
aud[1290]=16'he165;
aud[1291]=16'hc000;
aud[1292]=16'hac61;
aud[1293]=16'hb19e;
aud[1294]=16'hd0b0;
aud[1295]=16'h0;
aud[1296]=16'h2f50;
aud[1297]=16'h4e62;
aud[1298]=16'h539f;
aud[1299]=16'h4000;
aud[1300]=16'h1e9b;
aud[1301]=16'h0;
aud[1302]=16'hf352;
aud[1303]=16'h0;
aud[1304]=16'h22a3;
aud[1305]=16'h4e62;
aud[1306]=16'h723a;
aud[1307]=16'h7fff;
aud[1308]=16'h723a;
aud[1309]=16'h4e62;
aud[1310]=16'h22a3;
aud[1311]=16'h0;
aud[1312]=16'hf352;
aud[1313]=16'h0;
aud[1314]=16'h1e9b;
aud[1315]=16'h4000;
aud[1316]=16'h539f;
aud[1317]=16'h4e62;
aud[1318]=16'h2f50;
aud[1319]=16'h0;
aud[1320]=16'hd0b0;
aud[1321]=16'hb19e;
aud[1322]=16'hac61;
aud[1323]=16'hc000;
aud[1324]=16'he165;
aud[1325]=16'h0;
aud[1326]=16'hcae;
aud[1327]=16'h0;
aud[1328]=16'hdd5d;
aud[1329]=16'hb19e;
aud[1330]=16'h8dc6;
aud[1331]=16'h8000;
aud[1332]=16'h8dc6;
aud[1333]=16'hb19e;
aud[1334]=16'hdd5d;
aud[1335]=16'h0;
aud[1336]=16'hcae;
aud[1337]=16'h0;
aud[1338]=16'he165;
aud[1339]=16'hc000;
aud[1340]=16'hac61;
aud[1341]=16'hb19e;
aud[1342]=16'hd0b0;
aud[1343]=16'h0;
aud[1344]=16'h2f50;
aud[1345]=16'h4e62;
aud[1346]=16'h539f;
aud[1347]=16'h4000;
aud[1348]=16'h1e9b;
aud[1349]=16'h0;
aud[1350]=16'hf352;
aud[1351]=16'h0;
aud[1352]=16'h22a3;
aud[1353]=16'h4e62;
aud[1354]=16'h723a;
aud[1355]=16'h7fff;
aud[1356]=16'h723a;
aud[1357]=16'h4e62;
aud[1358]=16'h22a3;
aud[1359]=16'h0;
aud[1360]=16'hf352;
aud[1361]=16'h0;
aud[1362]=16'h1e9b;
aud[1363]=16'h4000;
aud[1364]=16'h539f;
aud[1365]=16'h4e62;
aud[1366]=16'h2f50;
aud[1367]=16'h0;
aud[1368]=16'hd0b0;
aud[1369]=16'hb19e;
aud[1370]=16'hac61;
aud[1371]=16'hc000;
aud[1372]=16'he165;
aud[1373]=16'h0;
aud[1374]=16'hcae;
aud[1375]=16'h0;
aud[1376]=16'hdd5d;
aud[1377]=16'hb19e;
aud[1378]=16'h8dc6;
aud[1379]=16'h8000;
aud[1380]=16'h8dc6;
aud[1381]=16'hb19e;
aud[1382]=16'hdd5d;
aud[1383]=16'h0;
aud[1384]=16'hcae;
aud[1385]=16'h0;
aud[1386]=16'he165;
aud[1387]=16'hc000;
aud[1388]=16'hac61;
aud[1389]=16'hb19e;
aud[1390]=16'hd0b0;
aud[1391]=16'h0;
aud[1392]=16'h2f50;
aud[1393]=16'h4e62;
aud[1394]=16'h539f;
aud[1395]=16'h4000;
aud[1396]=16'h1e9b;
aud[1397]=16'h0;
aud[1398]=16'hf352;
aud[1399]=16'h0;
aud[1400]=16'h22a3;
aud[1401]=16'h4e62;
aud[1402]=16'h723a;
aud[1403]=16'h7fff;
aud[1404]=16'h723a;
aud[1405]=16'h4e62;
aud[1406]=16'h22a3;
aud[1407]=16'h0;
aud[1408]=16'hf352;
aud[1409]=16'h0;
aud[1410]=16'h1e9b;
aud[1411]=16'h4000;
aud[1412]=16'h539f;
aud[1413]=16'h4e62;
aud[1414]=16'h2f50;
aud[1415]=16'h0;
aud[1416]=16'hd0b0;
aud[1417]=16'hb19e;
aud[1418]=16'hac61;
aud[1419]=16'hc000;
aud[1420]=16'he165;
aud[1421]=16'h0;
aud[1422]=16'hcae;
aud[1423]=16'h0;
aud[1424]=16'hdd5d;
aud[1425]=16'hb19e;
aud[1426]=16'h8dc6;
aud[1427]=16'h8000;
aud[1428]=16'h8dc6;
aud[1429]=16'hb19e;
aud[1430]=16'hdd5d;
aud[1431]=16'h0;
aud[1432]=16'hcae;
aud[1433]=16'h0;
aud[1434]=16'he165;
aud[1435]=16'hc000;
aud[1436]=16'hac61;
aud[1437]=16'hb19e;
aud[1438]=16'hd0b0;
aud[1439]=16'h0;
aud[1440]=16'h2f50;
aud[1441]=16'h4e62;
aud[1442]=16'h539f;
aud[1443]=16'h4000;
aud[1444]=16'h1e9b;
aud[1445]=16'h0;
aud[1446]=16'hf352;
aud[1447]=16'h0;
aud[1448]=16'h22a3;
aud[1449]=16'h4e62;
aud[1450]=16'h723a;
aud[1451]=16'h7fff;
aud[1452]=16'h723a;
aud[1453]=16'h4e62;
aud[1454]=16'h22a3;
aud[1455]=16'h0;
aud[1456]=16'hf352;
aud[1457]=16'h0;
aud[1458]=16'h1e9b;
aud[1459]=16'h4000;
aud[1460]=16'h539f;
aud[1461]=16'h4e62;
aud[1462]=16'h2f50;
aud[1463]=16'h0;
aud[1464]=16'hd0b0;
aud[1465]=16'hb19e;
aud[1466]=16'hac61;
aud[1467]=16'hc000;
aud[1468]=16'he165;
aud[1469]=16'h0;
aud[1470]=16'hcae;
aud[1471]=16'h0;
aud[1472]=16'hdd5d;
aud[1473]=16'hb19e;
aud[1474]=16'h8dc6;
aud[1475]=16'h8000;
aud[1476]=16'h8dc6;
aud[1477]=16'hb19e;
aud[1478]=16'hdd5d;
aud[1479]=16'h0;
aud[1480]=16'hcae;
aud[1481]=16'h0;
aud[1482]=16'he165;
aud[1483]=16'hc000;
aud[1484]=16'hac61;
aud[1485]=16'hb19e;
aud[1486]=16'hd0b0;
aud[1487]=16'h0;
aud[1488]=16'h2f50;
aud[1489]=16'h4e62;
aud[1490]=16'h539f;
aud[1491]=16'h4000;
aud[1492]=16'h1e9b;
aud[1493]=16'h0;
aud[1494]=16'hf352;
aud[1495]=16'h0;
aud[1496]=16'h22a3;
aud[1497]=16'h4e62;
aud[1498]=16'h723a;
aud[1499]=16'h7fff;
aud[1500]=16'h723a;
aud[1501]=16'h4e62;
aud[1502]=16'h22a3;
aud[1503]=16'h0;
aud[1504]=16'hf352;
aud[1505]=16'h0;
aud[1506]=16'h1e9b;
aud[1507]=16'h4000;
aud[1508]=16'h539f;
aud[1509]=16'h4e62;
aud[1510]=16'h2f50;
aud[1511]=16'h0;
aud[1512]=16'hd0b0;
aud[1513]=16'hb19e;
aud[1514]=16'hac61;
aud[1515]=16'hc000;
aud[1516]=16'he165;
aud[1517]=16'h0;
aud[1518]=16'hcae;
aud[1519]=16'h0;
aud[1520]=16'hdd5d;
aud[1521]=16'hb19e;
aud[1522]=16'h8dc6;
aud[1523]=16'h8000;
aud[1524]=16'h8dc6;
aud[1525]=16'hb19e;
aud[1526]=16'hdd5d;
aud[1527]=16'h0;
aud[1528]=16'hcae;
aud[1529]=16'h0;
aud[1530]=16'he165;
aud[1531]=16'hc000;
aud[1532]=16'hac61;
aud[1533]=16'hb19e;
aud[1534]=16'hd0b0;
aud[1535]=16'h0;
aud[1536]=16'h2f50;
aud[1537]=16'h4e62;
aud[1538]=16'h539f;
aud[1539]=16'h4000;
aud[1540]=16'h1e9b;
aud[1541]=16'h0;
aud[1542]=16'hf352;
aud[1543]=16'h0;
aud[1544]=16'h22a3;
aud[1545]=16'h4e62;
aud[1546]=16'h723a;
aud[1547]=16'h7fff;
aud[1548]=16'h723a;
aud[1549]=16'h4e62;
aud[1550]=16'h22a3;
aud[1551]=16'h0;
aud[1552]=16'hf352;
aud[1553]=16'h0;
aud[1554]=16'h1e9b;
aud[1555]=16'h4000;
aud[1556]=16'h539f;
aud[1557]=16'h4e62;
aud[1558]=16'h2f50;
aud[1559]=16'h0;
aud[1560]=16'hd0b0;
aud[1561]=16'hb19e;
aud[1562]=16'hac61;
aud[1563]=16'hc000;
aud[1564]=16'he165;
aud[1565]=16'h0;
aud[1566]=16'hcae;
aud[1567]=16'h0;
aud[1568]=16'hdd5d;
aud[1569]=16'hb19e;
aud[1570]=16'h8dc6;
aud[1571]=16'h8000;
aud[1572]=16'h8dc6;
aud[1573]=16'hb19e;
aud[1574]=16'hdd5d;
aud[1575]=16'h0;
aud[1576]=16'hcae;
aud[1577]=16'h0;
aud[1578]=16'he165;
aud[1579]=16'hc000;
aud[1580]=16'hac61;
aud[1581]=16'hb19e;
aud[1582]=16'hd0b0;
aud[1583]=16'h0;
aud[1584]=16'h2f50;
aud[1585]=16'h4e62;
aud[1586]=16'h539f;
aud[1587]=16'h4000;
aud[1588]=16'h1e9b;
aud[1589]=16'h0;
aud[1590]=16'hf352;
aud[1591]=16'h0;
aud[1592]=16'h22a3;
aud[1593]=16'h4e62;
aud[1594]=16'h723a;
aud[1595]=16'h7fff;
aud[1596]=16'h723a;
aud[1597]=16'h4e62;
aud[1598]=16'h22a3;
aud[1599]=16'h0;
aud[1600]=16'hf352;
aud[1601]=16'h0;
aud[1602]=16'h1e9b;
aud[1603]=16'h4000;
aud[1604]=16'h539f;
aud[1605]=16'h4e62;
aud[1606]=16'h2f50;
aud[1607]=16'h0;
aud[1608]=16'hd0b0;
aud[1609]=16'hb19e;
aud[1610]=16'hac61;
aud[1611]=16'hc000;
aud[1612]=16'he165;
aud[1613]=16'h0;
aud[1614]=16'hcae;
aud[1615]=16'h0;
aud[1616]=16'hdd5d;
aud[1617]=16'hb19e;
aud[1618]=16'h8dc6;
aud[1619]=16'h8000;
aud[1620]=16'h8dc6;
aud[1621]=16'hb19e;
aud[1622]=16'hdd5d;
aud[1623]=16'h0;
aud[1624]=16'hcae;
aud[1625]=16'h0;
aud[1626]=16'he165;
aud[1627]=16'hc000;
aud[1628]=16'hac61;
aud[1629]=16'hb19e;
aud[1630]=16'hd0b0;
aud[1631]=16'h0;
aud[1632]=16'h2f50;
aud[1633]=16'h4e62;
aud[1634]=16'h539f;
aud[1635]=16'h4000;
aud[1636]=16'h1e9b;
aud[1637]=16'h0;
aud[1638]=16'hf352;
aud[1639]=16'h0;
aud[1640]=16'h22a3;
aud[1641]=16'h4e62;
aud[1642]=16'h723a;
aud[1643]=16'h7fff;
aud[1644]=16'h723a;
aud[1645]=16'h4e62;
aud[1646]=16'h22a3;
aud[1647]=16'h0;
aud[1648]=16'hf352;
aud[1649]=16'h0;
aud[1650]=16'h1e9b;
aud[1651]=16'h4000;
aud[1652]=16'h539f;
aud[1653]=16'h4e62;
aud[1654]=16'h2f50;
aud[1655]=16'h0;
aud[1656]=16'hd0b0;
aud[1657]=16'hb19e;
aud[1658]=16'hac61;
aud[1659]=16'hc000;
aud[1660]=16'he165;
aud[1661]=16'h0;
aud[1662]=16'hcae;
aud[1663]=16'h0;
aud[1664]=16'hdd5d;
aud[1665]=16'hb19e;
aud[1666]=16'h8dc6;
aud[1667]=16'h8000;
aud[1668]=16'h8dc6;
aud[1669]=16'hb19e;
aud[1670]=16'hdd5d;
aud[1671]=16'h0;
aud[1672]=16'hcae;
aud[1673]=16'h0;
aud[1674]=16'he165;
aud[1675]=16'hc000;
aud[1676]=16'hac61;
aud[1677]=16'hb19e;
aud[1678]=16'hd0b0;
aud[1679]=16'h0;
aud[1680]=16'h2f50;
aud[1681]=16'h4e62;
aud[1682]=16'h539f;
aud[1683]=16'h4000;
aud[1684]=16'h1e9b;
aud[1685]=16'h0;
aud[1686]=16'hf352;
aud[1687]=16'h0;
aud[1688]=16'h22a3;
aud[1689]=16'h4e62;
aud[1690]=16'h723a;
aud[1691]=16'h7fff;
aud[1692]=16'h723a;
aud[1693]=16'h4e62;
aud[1694]=16'h22a3;
aud[1695]=16'h0;
aud[1696]=16'hf352;
aud[1697]=16'h0;
aud[1698]=16'h1e9b;
aud[1699]=16'h4000;
aud[1700]=16'h539f;
aud[1701]=16'h4e62;
aud[1702]=16'h2f50;
aud[1703]=16'h0;
aud[1704]=16'hd0b0;
aud[1705]=16'hb19e;
aud[1706]=16'hac61;
aud[1707]=16'hc000;
aud[1708]=16'he165;
aud[1709]=16'h0;
aud[1710]=16'hcae;
aud[1711]=16'h0;
aud[1712]=16'hdd5d;
aud[1713]=16'hb19e;
aud[1714]=16'h8dc6;
aud[1715]=16'h8000;
aud[1716]=16'h8dc6;
aud[1717]=16'hb19e;
aud[1718]=16'hdd5d;
aud[1719]=16'h0;
aud[1720]=16'hcae;
aud[1721]=16'h0;
aud[1722]=16'he165;
aud[1723]=16'hc000;
aud[1724]=16'hac61;
aud[1725]=16'hb19e;
aud[1726]=16'hd0b0;
aud[1727]=16'h0;
aud[1728]=16'h2f50;
aud[1729]=16'h4e62;
aud[1730]=16'h539f;
aud[1731]=16'h4000;
aud[1732]=16'h1e9b;
aud[1733]=16'h0;
aud[1734]=16'hf352;
aud[1735]=16'h0;
aud[1736]=16'h22a3;
aud[1737]=16'h4e62;
aud[1738]=16'h723a;
aud[1739]=16'h7fff;
aud[1740]=16'h723a;
aud[1741]=16'h4e62;
aud[1742]=16'h22a3;
aud[1743]=16'h0;
aud[1744]=16'hf352;
aud[1745]=16'h0;
aud[1746]=16'h1e9b;
aud[1747]=16'h4000;
aud[1748]=16'h539f;
aud[1749]=16'h4e62;
aud[1750]=16'h2f50;
aud[1751]=16'h0;
aud[1752]=16'hd0b0;
aud[1753]=16'hb19e;
aud[1754]=16'hac61;
aud[1755]=16'hc000;
aud[1756]=16'he165;
aud[1757]=16'h0;
aud[1758]=16'hcae;
aud[1759]=16'h0;
aud[1760]=16'hdd5d;
aud[1761]=16'hb19e;
aud[1762]=16'h8dc6;
aud[1763]=16'h8000;
aud[1764]=16'h8dc6;
aud[1765]=16'hb19e;
aud[1766]=16'hdd5d;
aud[1767]=16'h0;
aud[1768]=16'hcae;
aud[1769]=16'h0;
aud[1770]=16'he165;
aud[1771]=16'hc000;
aud[1772]=16'hac61;
aud[1773]=16'hb19e;
aud[1774]=16'hd0b0;
aud[1775]=16'h0;
aud[1776]=16'h2f50;
aud[1777]=16'h4e62;
aud[1778]=16'h539f;
aud[1779]=16'h4000;
aud[1780]=16'h1e9b;
aud[1781]=16'h0;
aud[1782]=16'hf352;
aud[1783]=16'h0;
aud[1784]=16'h22a3;
aud[1785]=16'h4e62;
aud[1786]=16'h723a;
aud[1787]=16'h7fff;
aud[1788]=16'h723a;
aud[1789]=16'h4e62;
aud[1790]=16'h22a3;
aud[1791]=16'h0;
aud[1792]=16'hf352;
aud[1793]=16'h0;
aud[1794]=16'h1e9b;
aud[1795]=16'h4000;
aud[1796]=16'h539f;
aud[1797]=16'h4e62;
aud[1798]=16'h2f50;
aud[1799]=16'h0;
aud[1800]=16'hd0b0;
aud[1801]=16'hb19e;
aud[1802]=16'hac61;
aud[1803]=16'hc000;
aud[1804]=16'he165;
aud[1805]=16'h0;
aud[1806]=16'hcae;
aud[1807]=16'h0;
aud[1808]=16'hdd5d;
aud[1809]=16'hb19e;
aud[1810]=16'h8dc6;
aud[1811]=16'h8000;
aud[1812]=16'h8dc6;
aud[1813]=16'hb19e;
aud[1814]=16'hdd5d;
aud[1815]=16'h0;
aud[1816]=16'hcae;
aud[1817]=16'h0;
aud[1818]=16'he165;
aud[1819]=16'hc000;
aud[1820]=16'hac61;
aud[1821]=16'hb19e;
aud[1822]=16'hd0b0;
aud[1823]=16'h0;
aud[1824]=16'h2f50;
aud[1825]=16'h4e62;
aud[1826]=16'h539f;
aud[1827]=16'h4000;
aud[1828]=16'h1e9b;
aud[1829]=16'h0;
aud[1830]=16'hf352;
aud[1831]=16'h0;
aud[1832]=16'h22a3;
aud[1833]=16'h4e62;
aud[1834]=16'h723a;
aud[1835]=16'h7fff;
aud[1836]=16'h723a;
aud[1837]=16'h4e62;
aud[1838]=16'h22a3;
aud[1839]=16'h0;
aud[1840]=16'hf352;
aud[1841]=16'h0;
aud[1842]=16'h1e9b;
aud[1843]=16'h4000;
aud[1844]=16'h539f;
aud[1845]=16'h4e62;
aud[1846]=16'h2f50;
aud[1847]=16'h0;
aud[1848]=16'hd0b0;
aud[1849]=16'hb19e;
aud[1850]=16'hac61;
aud[1851]=16'hc000;
aud[1852]=16'he165;
aud[1853]=16'h0;
aud[1854]=16'hcae;
aud[1855]=16'h0;
aud[1856]=16'hdd5d;
aud[1857]=16'hb19e;
aud[1858]=16'h8dc6;
aud[1859]=16'h8000;
aud[1860]=16'h8dc6;
aud[1861]=16'hb19e;
aud[1862]=16'hdd5d;
aud[1863]=16'h0;
aud[1864]=16'hcae;
aud[1865]=16'h0;
aud[1866]=16'he165;
aud[1867]=16'hc000;
aud[1868]=16'hac61;
aud[1869]=16'hb19e;
aud[1870]=16'hd0b0;
aud[1871]=16'h0;
aud[1872]=16'h2f50;
aud[1873]=16'h4e62;
aud[1874]=16'h539f;
aud[1875]=16'h4000;
aud[1876]=16'h1e9b;
aud[1877]=16'h0;
aud[1878]=16'hf352;
aud[1879]=16'h0;
aud[1880]=16'h22a3;
aud[1881]=16'h4e62;
aud[1882]=16'h723a;
aud[1883]=16'h7fff;
aud[1884]=16'h723a;
aud[1885]=16'h4e62;
aud[1886]=16'h22a3;
aud[1887]=16'h0;
aud[1888]=16'hf352;
aud[1889]=16'h0;
aud[1890]=16'h1e9b;
aud[1891]=16'h4000;
aud[1892]=16'h539f;
aud[1893]=16'h4e62;
aud[1894]=16'h2f50;
aud[1895]=16'h0;
aud[1896]=16'hd0b0;
aud[1897]=16'hb19e;
aud[1898]=16'hac61;
aud[1899]=16'hc000;
aud[1900]=16'he165;
aud[1901]=16'h0;
aud[1902]=16'hcae;
aud[1903]=16'h0;
aud[1904]=16'hdd5d;
aud[1905]=16'hb19e;
aud[1906]=16'h8dc6;
aud[1907]=16'h8000;
aud[1908]=16'h8dc6;
aud[1909]=16'hb19e;
aud[1910]=16'hdd5d;
aud[1911]=16'h0;
aud[1912]=16'hcae;
aud[1913]=16'h0;
aud[1914]=16'he165;
aud[1915]=16'hc000;
aud[1916]=16'hac61;
aud[1917]=16'hb19e;
aud[1918]=16'hd0b0;
aud[1919]=16'h0;
aud[1920]=16'h2f50;
aud[1921]=16'h4e62;
aud[1922]=16'h539f;
aud[1923]=16'h4000;
aud[1924]=16'h1e9b;
aud[1925]=16'h0;
aud[1926]=16'hf352;
aud[1927]=16'h0;
aud[1928]=16'h22a3;
aud[1929]=16'h4e62;
aud[1930]=16'h723a;
aud[1931]=16'h7fff;
aud[1932]=16'h723a;
aud[1933]=16'h4e62;
aud[1934]=16'h22a3;
aud[1935]=16'h0;
aud[1936]=16'hf352;
aud[1937]=16'h0;
aud[1938]=16'h1e9b;
aud[1939]=16'h4000;
aud[1940]=16'h539f;
aud[1941]=16'h4e62;
aud[1942]=16'h2f50;
aud[1943]=16'h0;
aud[1944]=16'hd0b0;
aud[1945]=16'hb19e;
aud[1946]=16'hac61;
aud[1947]=16'hc000;
aud[1948]=16'he165;
aud[1949]=16'h0;
aud[1950]=16'hcae;
aud[1951]=16'h0;
aud[1952]=16'hdd5d;
aud[1953]=16'hb19e;
aud[1954]=16'h8dc6;
aud[1955]=16'h8000;
aud[1956]=16'h8dc6;
aud[1957]=16'hb19e;
aud[1958]=16'hdd5d;
aud[1959]=16'h0;
aud[1960]=16'hcae;
aud[1961]=16'h0;
aud[1962]=16'he165;
aud[1963]=16'hc000;
aud[1964]=16'hac61;
aud[1965]=16'hb19e;
aud[1966]=16'hd0b0;
aud[1967]=16'h0;
aud[1968]=16'h2f50;
aud[1969]=16'h4e62;
aud[1970]=16'h539f;
aud[1971]=16'h4000;
aud[1972]=16'h1e9b;
aud[1973]=16'h0;
aud[1974]=16'hf352;
aud[1975]=16'h0;
aud[1976]=16'h22a3;
aud[1977]=16'h4e62;
aud[1978]=16'h723a;
aud[1979]=16'h7fff;
aud[1980]=16'h723a;
aud[1981]=16'h4e62;
aud[1982]=16'h22a3;
aud[1983]=16'h0;
aud[1984]=16'hf352;
aud[1985]=16'h0;
aud[1986]=16'h1e9b;
aud[1987]=16'h4000;
aud[1988]=16'h539f;
aud[1989]=16'h4e62;
aud[1990]=16'h2f50;
aud[1991]=16'h0;
aud[1992]=16'hd0b0;
aud[1993]=16'hb19e;
aud[1994]=16'hac61;
aud[1995]=16'hc000;
aud[1996]=16'he165;
aud[1997]=16'h0;
aud[1998]=16'hcae;
aud[1999]=16'h0;

end


endmodule