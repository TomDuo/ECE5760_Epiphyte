//=============================================================================
// Lab 1 - Cellular Automata Control File
//
// Authors:
//  Connor Archard
//  Kevin Kreher
//  Noah Levy
//
// Date:
//  Feb 3, 2016
//=============================================================================

module lab1_ctrl(
	input clk,
	input SW[17:0]),
	
	
	assign f=(x1 & x2);
endmodule