module testVect (
output reg signed [15:0] aud [0:49999]
);

initial begin
aud[0]=16'h15;
aud[1]=16'h2b;
aud[2]=16'h40;
aud[3]=16'h56;
aud[4]=16'h6b;
aud[5]=16'h81;
aud[6]=16'h96;
aud[7]=16'hac;
aud[8]=16'hc1;
aud[9]=16'hd6;
aud[10]=16'hec;
aud[11]=16'h101;
aud[12]=16'h117;
aud[13]=16'h12c;
aud[14]=16'h142;
aud[15]=16'h157;
aud[16]=16'h16d;
aud[17]=16'h182;
aud[18]=16'h197;
aud[19]=16'h1ad;
aud[20]=16'h1c2;
aud[21]=16'h1d8;
aud[22]=16'h1ed;
aud[23]=16'h203;
aud[24]=16'h218;
aud[25]=16'h22e;
aud[26]=16'h243;
aud[27]=16'h258;
aud[28]=16'h26e;
aud[29]=16'h283;
aud[30]=16'h299;
aud[31]=16'h2ae;
aud[32]=16'h2c4;
aud[33]=16'h2d9;
aud[34]=16'h2ee;
aud[35]=16'h304;
aud[36]=16'h319;
aud[37]=16'h32f;
aud[38]=16'h344;
aud[39]=16'h359;
aud[40]=16'h36f;
aud[41]=16'h384;
aud[42]=16'h39a;
aud[43]=16'h3af;
aud[44]=16'h3c5;
aud[45]=16'h3da;
aud[46]=16'h3ef;
aud[47]=16'h405;
aud[48]=16'h41a;
aud[49]=16'h430;
aud[50]=16'h445;
aud[51]=16'h45a;
aud[52]=16'h470;
aud[53]=16'h485;
aud[54]=16'h49b;
aud[55]=16'h4b0;
aud[56]=16'h4c5;
aud[57]=16'h4db;
aud[58]=16'h4f0;
aud[59]=16'h505;
aud[60]=16'h51b;
aud[61]=16'h530;
aud[62]=16'h546;
aud[63]=16'h55b;
aud[64]=16'h570;
aud[65]=16'h586;
aud[66]=16'h59b;
aud[67]=16'h5b0;
aud[68]=16'h5c6;
aud[69]=16'h5db;
aud[70]=16'h5f1;
aud[71]=16'h606;
aud[72]=16'h61b;
aud[73]=16'h631;
aud[74]=16'h646;
aud[75]=16'h65b;
aud[76]=16'h671;
aud[77]=16'h686;
aud[78]=16'h69b;
aud[79]=16'h6b1;
aud[80]=16'h6c6;
aud[81]=16'h6db;
aud[82]=16'h6f1;
aud[83]=16'h706;
aud[84]=16'h71b;
aud[85]=16'h731;
aud[86]=16'h746;
aud[87]=16'h75b;
aud[88]=16'h770;
aud[89]=16'h786;
aud[90]=16'h79b;
aud[91]=16'h7b0;
aud[92]=16'h7c6;
aud[93]=16'h7db;
aud[94]=16'h7f0;
aud[95]=16'h805;
aud[96]=16'h81b;
aud[97]=16'h830;
aud[98]=16'h845;
aud[99]=16'h85b;
aud[100]=16'h870;
aud[101]=16'h885;
aud[102]=16'h89a;
aud[103]=16'h8b0;
aud[104]=16'h8c5;
aud[105]=16'h8da;
aud[106]=16'h8ef;
aud[107]=16'h905;
aud[108]=16'h91a;
aud[109]=16'h92f;
aud[110]=16'h944;
aud[111]=16'h959;
aud[112]=16'h96f;
aud[113]=16'h984;
aud[114]=16'h999;
aud[115]=16'h9ae;
aud[116]=16'h9c3;
aud[117]=16'h9d9;
aud[118]=16'h9ee;
aud[119]=16'ha03;
aud[120]=16'ha18;
aud[121]=16'ha2d;
aud[122]=16'ha43;
aud[123]=16'ha58;
aud[124]=16'ha6d;
aud[125]=16'ha82;
aud[126]=16'ha97;
aud[127]=16'haac;
aud[128]=16'hac1;
aud[129]=16'had7;
aud[130]=16'haec;
aud[131]=16'hb01;
aud[132]=16'hb16;
aud[133]=16'hb2b;
aud[134]=16'hb40;
aud[135]=16'hb55;
aud[136]=16'hb6a;
aud[137]=16'hb80;
aud[138]=16'hb95;
aud[139]=16'hbaa;
aud[140]=16'hbbf;
aud[141]=16'hbd4;
aud[142]=16'hbe9;
aud[143]=16'hbfe;
aud[144]=16'hc13;
aud[145]=16'hc28;
aud[146]=16'hc3d;
aud[147]=16'hc52;
aud[148]=16'hc67;
aud[149]=16'hc7c;
aud[150]=16'hc91;
aud[151]=16'hca6;
aud[152]=16'hcbb;
aud[153]=16'hcd0;
aud[154]=16'hce5;
aud[155]=16'hcfa;
aud[156]=16'hd0f;
aud[157]=16'hd24;
aud[158]=16'hd39;
aud[159]=16'hd4e;
aud[160]=16'hd63;
aud[161]=16'hd78;
aud[162]=16'hd8d;
aud[163]=16'hda2;
aud[164]=16'hdb7;
aud[165]=16'hdcc;
aud[166]=16'hde1;
aud[167]=16'hdf6;
aud[168]=16'he0b;
aud[169]=16'he20;
aud[170]=16'he35;
aud[171]=16'he4a;
aud[172]=16'he5f;
aud[173]=16'he74;
aud[174]=16'he88;
aud[175]=16'he9d;
aud[176]=16'heb2;
aud[177]=16'hec7;
aud[178]=16'hedc;
aud[179]=16'hef1;
aud[180]=16'hf06;
aud[181]=16'hf1a;
aud[182]=16'hf2f;
aud[183]=16'hf44;
aud[184]=16'hf59;
aud[185]=16'hf6e;
aud[186]=16'hf83;
aud[187]=16'hf97;
aud[188]=16'hfac;
aud[189]=16'hfc1;
aud[190]=16'hfd6;
aud[191]=16'hfeb;
aud[192]=16'hfff;
aud[193]=16'h1014;
aud[194]=16'h1029;
aud[195]=16'h103e;
aud[196]=16'h1052;
aud[197]=16'h1067;
aud[198]=16'h107c;
aud[199]=16'h1090;
aud[200]=16'h10a5;
aud[201]=16'h10ba;
aud[202]=16'h10cf;
aud[203]=16'h10e3;
aud[204]=16'h10f8;
aud[205]=16'h110d;
aud[206]=16'h1121;
aud[207]=16'h1136;
aud[208]=16'h114b;
aud[209]=16'h115f;
aud[210]=16'h1174;
aud[211]=16'h1189;
aud[212]=16'h119d;
aud[213]=16'h11b2;
aud[214]=16'h11c6;
aud[215]=16'h11db;
aud[216]=16'h11f0;
aud[217]=16'h1204;
aud[218]=16'h1219;
aud[219]=16'h122d;
aud[220]=16'h1242;
aud[221]=16'h1256;
aud[222]=16'h126b;
aud[223]=16'h127f;
aud[224]=16'h1294;
aud[225]=16'h12a9;
aud[226]=16'h12bd;
aud[227]=16'h12d2;
aud[228]=16'h12e6;
aud[229]=16'h12fb;
aud[230]=16'h130f;
aud[231]=16'h1323;
aud[232]=16'h1338;
aud[233]=16'h134c;
aud[234]=16'h1361;
aud[235]=16'h1375;
aud[236]=16'h138a;
aud[237]=16'h139e;
aud[238]=16'h13b3;
aud[239]=16'h13c7;
aud[240]=16'h13db;
aud[241]=16'h13f0;
aud[242]=16'h1404;
aud[243]=16'h1418;
aud[244]=16'h142d;
aud[245]=16'h1441;
aud[246]=16'h1455;
aud[247]=16'h146a;
aud[248]=16'h147e;
aud[249]=16'h1492;
aud[250]=16'h14a7;
aud[251]=16'h14bb;
aud[252]=16'h14cf;
aud[253]=16'h14e4;
aud[254]=16'h14f8;
aud[255]=16'h150c;
aud[256]=16'h1520;
aud[257]=16'h1535;
aud[258]=16'h1549;
aud[259]=16'h155d;
aud[260]=16'h1571;
aud[261]=16'h1586;
aud[262]=16'h159a;
aud[263]=16'h15ae;
aud[264]=16'h15c2;
aud[265]=16'h15d6;
aud[266]=16'h15ea;
aud[267]=16'h15ff;
aud[268]=16'h1613;
aud[269]=16'h1627;
aud[270]=16'h163b;
aud[271]=16'h164f;
aud[272]=16'h1663;
aud[273]=16'h1677;
aud[274]=16'h168b;
aud[275]=16'h169f;
aud[276]=16'h16b3;
aud[277]=16'h16c7;
aud[278]=16'h16db;
aud[279]=16'h16f0;
aud[280]=16'h1704;
aud[281]=16'h1718;
aud[282]=16'h172c;
aud[283]=16'h1740;
aud[284]=16'h1753;
aud[285]=16'h1767;
aud[286]=16'h177b;
aud[287]=16'h178f;
aud[288]=16'h17a3;
aud[289]=16'h17b7;
aud[290]=16'h17cb;
aud[291]=16'h17df;
aud[292]=16'h17f3;
aud[293]=16'h1807;
aud[294]=16'h181b;
aud[295]=16'h182f;
aud[296]=16'h1842;
aud[297]=16'h1856;
aud[298]=16'h186a;
aud[299]=16'h187e;
aud[300]=16'h1892;
aud[301]=16'h18a5;
aud[302]=16'h18b9;
aud[303]=16'h18cd;
aud[304]=16'h18e1;
aud[305]=16'h18f5;
aud[306]=16'h1908;
aud[307]=16'h191c;
aud[308]=16'h1930;
aud[309]=16'h1943;
aud[310]=16'h1957;
aud[311]=16'h196b;
aud[312]=16'h197f;
aud[313]=16'h1992;
aud[314]=16'h19a6;
aud[315]=16'h19ba;
aud[316]=16'h19cd;
aud[317]=16'h19e1;
aud[318]=16'h19f4;
aud[319]=16'h1a08;
aud[320]=16'h1a1c;
aud[321]=16'h1a2f;
aud[322]=16'h1a43;
aud[323]=16'h1a56;
aud[324]=16'h1a6a;
aud[325]=16'h1a7d;
aud[326]=16'h1a91;
aud[327]=16'h1aa4;
aud[328]=16'h1ab8;
aud[329]=16'h1acb;
aud[330]=16'h1adf;
aud[331]=16'h1af2;
aud[332]=16'h1b06;
aud[333]=16'h1b19;
aud[334]=16'h1b2d;
aud[335]=16'h1b40;
aud[336]=16'h1b53;
aud[337]=16'h1b67;
aud[338]=16'h1b7a;
aud[339]=16'h1b8d;
aud[340]=16'h1ba1;
aud[341]=16'h1bb4;
aud[342]=16'h1bc8;
aud[343]=16'h1bdb;
aud[344]=16'h1bee;
aud[345]=16'h1c01;
aud[346]=16'h1c15;
aud[347]=16'h1c28;
aud[348]=16'h1c3b;
aud[349]=16'h1c4e;
aud[350]=16'h1c62;
aud[351]=16'h1c75;
aud[352]=16'h1c88;
aud[353]=16'h1c9b;
aud[354]=16'h1cae;
aud[355]=16'h1cc2;
aud[356]=16'h1cd5;
aud[357]=16'h1ce8;
aud[358]=16'h1cfb;
aud[359]=16'h1d0e;
aud[360]=16'h1d21;
aud[361]=16'h1d34;
aud[362]=16'h1d47;
aud[363]=16'h1d5b;
aud[364]=16'h1d6e;
aud[365]=16'h1d81;
aud[366]=16'h1d94;
aud[367]=16'h1da7;
aud[368]=16'h1dba;
aud[369]=16'h1dcd;
aud[370]=16'h1de0;
aud[371]=16'h1df3;
aud[372]=16'h1e06;
aud[373]=16'h1e18;
aud[374]=16'h1e2b;
aud[375]=16'h1e3e;
aud[376]=16'h1e51;
aud[377]=16'h1e64;
aud[378]=16'h1e77;
aud[379]=16'h1e8a;
aud[380]=16'h1e9d;
aud[381]=16'h1eaf;
aud[382]=16'h1ec2;
aud[383]=16'h1ed5;
aud[384]=16'h1ee8;
aud[385]=16'h1efb;
aud[386]=16'h1f0d;
aud[387]=16'h1f20;
aud[388]=16'h1f33;
aud[389]=16'h1f46;
aud[390]=16'h1f58;
aud[391]=16'h1f6b;
aud[392]=16'h1f7e;
aud[393]=16'h1f90;
aud[394]=16'h1fa3;
aud[395]=16'h1fb6;
aud[396]=16'h1fc8;
aud[397]=16'h1fdb;
aud[398]=16'h1fed;
aud[399]=16'h2000;
aud[400]=16'h2013;
aud[401]=16'h2025;
aud[402]=16'h2038;
aud[403]=16'h204a;
aud[404]=16'h205d;
aud[405]=16'h206f;
aud[406]=16'h2082;
aud[407]=16'h2094;
aud[408]=16'h20a7;
aud[409]=16'h20b9;
aud[410]=16'h20cb;
aud[411]=16'h20de;
aud[412]=16'h20f0;
aud[413]=16'h2103;
aud[414]=16'h2115;
aud[415]=16'h2127;
aud[416]=16'h213a;
aud[417]=16'h214c;
aud[418]=16'h215e;
aud[419]=16'h2171;
aud[420]=16'h2183;
aud[421]=16'h2195;
aud[422]=16'h21a7;
aud[423]=16'h21ba;
aud[424]=16'h21cc;
aud[425]=16'h21de;
aud[426]=16'h21f0;
aud[427]=16'h2202;
aud[428]=16'h2215;
aud[429]=16'h2227;
aud[430]=16'h2239;
aud[431]=16'h224b;
aud[432]=16'h225d;
aud[433]=16'h226f;
aud[434]=16'h2281;
aud[435]=16'h2293;
aud[436]=16'h22a5;
aud[437]=16'h22b7;
aud[438]=16'h22c9;
aud[439]=16'h22db;
aud[440]=16'h22ed;
aud[441]=16'h22ff;
aud[442]=16'h2311;
aud[443]=16'h2323;
aud[444]=16'h2335;
aud[445]=16'h2347;
aud[446]=16'h2359;
aud[447]=16'h236b;
aud[448]=16'h237d;
aud[449]=16'h238e;
aud[450]=16'h23a0;
aud[451]=16'h23b2;
aud[452]=16'h23c4;
aud[453]=16'h23d6;
aud[454]=16'h23e7;
aud[455]=16'h23f9;
aud[456]=16'h240b;
aud[457]=16'h241d;
aud[458]=16'h242e;
aud[459]=16'h2440;
aud[460]=16'h2452;
aud[461]=16'h2463;
aud[462]=16'h2475;
aud[463]=16'h2487;
aud[464]=16'h2498;
aud[465]=16'h24aa;
aud[466]=16'h24bb;
aud[467]=16'h24cd;
aud[468]=16'h24de;
aud[469]=16'h24f0;
aud[470]=16'h2501;
aud[471]=16'h2513;
aud[472]=16'h2524;
aud[473]=16'h2536;
aud[474]=16'h2547;
aud[475]=16'h2559;
aud[476]=16'h256a;
aud[477]=16'h257c;
aud[478]=16'h258d;
aud[479]=16'h259e;
aud[480]=16'h25b0;
aud[481]=16'h25c1;
aud[482]=16'h25d2;
aud[483]=16'h25e4;
aud[484]=16'h25f5;
aud[485]=16'h2606;
aud[486]=16'h2617;
aud[487]=16'h2629;
aud[488]=16'h263a;
aud[489]=16'h264b;
aud[490]=16'h265c;
aud[491]=16'h266d;
aud[492]=16'h267e;
aud[493]=16'h2690;
aud[494]=16'h26a1;
aud[495]=16'h26b2;
aud[496]=16'h26c3;
aud[497]=16'h26d4;
aud[498]=16'h26e5;
aud[499]=16'h26f6;
aud[500]=16'h2707;
aud[501]=16'h2718;
aud[502]=16'h2729;
aud[503]=16'h273a;
aud[504]=16'h274b;
aud[505]=16'h275c;
aud[506]=16'h276d;
aud[507]=16'h277e;
aud[508]=16'h278e;
aud[509]=16'h279f;
aud[510]=16'h27b0;
aud[511]=16'h27c1;
aud[512]=16'h27d2;
aud[513]=16'h27e2;
aud[514]=16'h27f3;
aud[515]=16'h2804;
aud[516]=16'h2815;
aud[517]=16'h2825;
aud[518]=16'h2836;
aud[519]=16'h2847;
aud[520]=16'h2857;
aud[521]=16'h2868;
aud[522]=16'h2879;
aud[523]=16'h2889;
aud[524]=16'h289a;
aud[525]=16'h28aa;
aud[526]=16'h28bb;
aud[527]=16'h28cc;
aud[528]=16'h28dc;
aud[529]=16'h28ed;
aud[530]=16'h28fd;
aud[531]=16'h290e;
aud[532]=16'h291e;
aud[533]=16'h292e;
aud[534]=16'h293f;
aud[535]=16'h294f;
aud[536]=16'h2960;
aud[537]=16'h2970;
aud[538]=16'h2980;
aud[539]=16'h2991;
aud[540]=16'h29a1;
aud[541]=16'h29b1;
aud[542]=16'h29c1;
aud[543]=16'h29d2;
aud[544]=16'h29e2;
aud[545]=16'h29f2;
aud[546]=16'h2a02;
aud[547]=16'h2a12;
aud[548]=16'h2a23;
aud[549]=16'h2a33;
aud[550]=16'h2a43;
aud[551]=16'h2a53;
aud[552]=16'h2a63;
aud[553]=16'h2a73;
aud[554]=16'h2a83;
aud[555]=16'h2a93;
aud[556]=16'h2aa3;
aud[557]=16'h2ab3;
aud[558]=16'h2ac3;
aud[559]=16'h2ad3;
aud[560]=16'h2ae3;
aud[561]=16'h2af3;
aud[562]=16'h2b03;
aud[563]=16'h2b13;
aud[564]=16'h2b22;
aud[565]=16'h2b32;
aud[566]=16'h2b42;
aud[567]=16'h2b52;
aud[568]=16'h2b62;
aud[569]=16'h2b71;
aud[570]=16'h2b81;
aud[571]=16'h2b91;
aud[572]=16'h2ba1;
aud[573]=16'h2bb0;
aud[574]=16'h2bc0;
aud[575]=16'h2bd0;
aud[576]=16'h2bdf;
aud[577]=16'h2bef;
aud[578]=16'h2bfe;
aud[579]=16'h2c0e;
aud[580]=16'h2c1e;
aud[581]=16'h2c2d;
aud[582]=16'h2c3d;
aud[583]=16'h2c4c;
aud[584]=16'h2c5c;
aud[585]=16'h2c6b;
aud[586]=16'h2c7a;
aud[587]=16'h2c8a;
aud[588]=16'h2c99;
aud[589]=16'h2ca9;
aud[590]=16'h2cb8;
aud[591]=16'h2cc7;
aud[592]=16'h2cd7;
aud[593]=16'h2ce6;
aud[594]=16'h2cf5;
aud[595]=16'h2d04;
aud[596]=16'h2d14;
aud[597]=16'h2d23;
aud[598]=16'h2d32;
aud[599]=16'h2d41;
aud[600]=16'h2d50;
aud[601]=16'h2d60;
aud[602]=16'h2d6f;
aud[603]=16'h2d7e;
aud[604]=16'h2d8d;
aud[605]=16'h2d9c;
aud[606]=16'h2dab;
aud[607]=16'h2dba;
aud[608]=16'h2dc9;
aud[609]=16'h2dd8;
aud[610]=16'h2de7;
aud[611]=16'h2df6;
aud[612]=16'h2e05;
aud[613]=16'h2e14;
aud[614]=16'h2e22;
aud[615]=16'h2e31;
aud[616]=16'h2e40;
aud[617]=16'h2e4f;
aud[618]=16'h2e5e;
aud[619]=16'h2e6d;
aud[620]=16'h2e7b;
aud[621]=16'h2e8a;
aud[622]=16'h2e99;
aud[623]=16'h2ea7;
aud[624]=16'h2eb6;
aud[625]=16'h2ec5;
aud[626]=16'h2ed3;
aud[627]=16'h2ee2;
aud[628]=16'h2ef1;
aud[629]=16'h2eff;
aud[630]=16'h2f0e;
aud[631]=16'h2f1c;
aud[632]=16'h2f2b;
aud[633]=16'h2f39;
aud[634]=16'h2f48;
aud[635]=16'h2f56;
aud[636]=16'h2f65;
aud[637]=16'h2f73;
aud[638]=16'h2f81;
aud[639]=16'h2f90;
aud[640]=16'h2f9e;
aud[641]=16'h2fac;
aud[642]=16'h2fbb;
aud[643]=16'h2fc9;
aud[644]=16'h2fd7;
aud[645]=16'h2fe5;
aud[646]=16'h2ff4;
aud[647]=16'h3002;
aud[648]=16'h3010;
aud[649]=16'h301e;
aud[650]=16'h302c;
aud[651]=16'h303a;
aud[652]=16'h3048;
aud[653]=16'h3057;
aud[654]=16'h3065;
aud[655]=16'h3073;
aud[656]=16'h3081;
aud[657]=16'h308f;
aud[658]=16'h309d;
aud[659]=16'h30aa;
aud[660]=16'h30b8;
aud[661]=16'h30c6;
aud[662]=16'h30d4;
aud[663]=16'h30e2;
aud[664]=16'h30f0;
aud[665]=16'h30fe;
aud[666]=16'h310b;
aud[667]=16'h3119;
aud[668]=16'h3127;
aud[669]=16'h3135;
aud[670]=16'h3142;
aud[671]=16'h3150;
aud[672]=16'h315e;
aud[673]=16'h316b;
aud[674]=16'h3179;
aud[675]=16'h3187;
aud[676]=16'h3194;
aud[677]=16'h31a2;
aud[678]=16'h31af;
aud[679]=16'h31bd;
aud[680]=16'h31ca;
aud[681]=16'h31d8;
aud[682]=16'h31e5;
aud[683]=16'h31f3;
aud[684]=16'h3200;
aud[685]=16'h320d;
aud[686]=16'h321b;
aud[687]=16'h3228;
aud[688]=16'h3235;
aud[689]=16'h3243;
aud[690]=16'h3250;
aud[691]=16'h325d;
aud[692]=16'h326a;
aud[693]=16'h3278;
aud[694]=16'h3285;
aud[695]=16'h3292;
aud[696]=16'h329f;
aud[697]=16'h32ac;
aud[698]=16'h32b9;
aud[699]=16'h32c6;
aud[700]=16'h32d3;
aud[701]=16'h32e0;
aud[702]=16'h32ed;
aud[703]=16'h32fa;
aud[704]=16'h3307;
aud[705]=16'h3314;
aud[706]=16'h3321;
aud[707]=16'h332e;
aud[708]=16'h333b;
aud[709]=16'h3348;
aud[710]=16'h3355;
aud[711]=16'h3361;
aud[712]=16'h336e;
aud[713]=16'h337b;
aud[714]=16'h3388;
aud[715]=16'h3394;
aud[716]=16'h33a1;
aud[717]=16'h33ae;
aud[718]=16'h33ba;
aud[719]=16'h33c7;
aud[720]=16'h33d4;
aud[721]=16'h33e0;
aud[722]=16'h33ed;
aud[723]=16'h33f9;
aud[724]=16'h3406;
aud[725]=16'h3412;
aud[726]=16'h341f;
aud[727]=16'h342b;
aud[728]=16'h3437;
aud[729]=16'h3444;
aud[730]=16'h3450;
aud[731]=16'h345d;
aud[732]=16'h3469;
aud[733]=16'h3475;
aud[734]=16'h3481;
aud[735]=16'h348e;
aud[736]=16'h349a;
aud[737]=16'h34a6;
aud[738]=16'h34b2;
aud[739]=16'h34be;
aud[740]=16'h34cb;
aud[741]=16'h34d7;
aud[742]=16'h34e3;
aud[743]=16'h34ef;
aud[744]=16'h34fb;
aud[745]=16'h3507;
aud[746]=16'h3513;
aud[747]=16'h351f;
aud[748]=16'h352b;
aud[749]=16'h3537;
aud[750]=16'h3543;
aud[751]=16'h354f;
aud[752]=16'h355a;
aud[753]=16'h3566;
aud[754]=16'h3572;
aud[755]=16'h357e;
aud[756]=16'h358a;
aud[757]=16'h3595;
aud[758]=16'h35a1;
aud[759]=16'h35ad;
aud[760]=16'h35b8;
aud[761]=16'h35c4;
aud[762]=16'h35d0;
aud[763]=16'h35db;
aud[764]=16'h35e7;
aud[765]=16'h35f2;
aud[766]=16'h35fe;
aud[767]=16'h3609;
aud[768]=16'h3615;
aud[769]=16'h3620;
aud[770]=16'h362c;
aud[771]=16'h3637;
aud[772]=16'h3643;
aud[773]=16'h364e;
aud[774]=16'h3659;
aud[775]=16'h3665;
aud[776]=16'h3670;
aud[777]=16'h367b;
aud[778]=16'h3686;
aud[779]=16'h3692;
aud[780]=16'h369d;
aud[781]=16'h36a8;
aud[782]=16'h36b3;
aud[783]=16'h36be;
aud[784]=16'h36c9;
aud[785]=16'h36d4;
aud[786]=16'h36e0;
aud[787]=16'h36eb;
aud[788]=16'h36f6;
aud[789]=16'h3701;
aud[790]=16'h370b;
aud[791]=16'h3716;
aud[792]=16'h3721;
aud[793]=16'h372c;
aud[794]=16'h3737;
aud[795]=16'h3742;
aud[796]=16'h374d;
aud[797]=16'h3757;
aud[798]=16'h3762;
aud[799]=16'h376d;
aud[800]=16'h3778;
aud[801]=16'h3782;
aud[802]=16'h378d;
aud[803]=16'h3798;
aud[804]=16'h37a2;
aud[805]=16'h37ad;
aud[806]=16'h37b7;
aud[807]=16'h37c2;
aud[808]=16'h37cc;
aud[809]=16'h37d7;
aud[810]=16'h37e1;
aud[811]=16'h37ec;
aud[812]=16'h37f6;
aud[813]=16'h3801;
aud[814]=16'h380b;
aud[815]=16'h3815;
aud[816]=16'h3820;
aud[817]=16'h382a;
aud[818]=16'h3834;
aud[819]=16'h383f;
aud[820]=16'h3849;
aud[821]=16'h3853;
aud[822]=16'h385d;
aud[823]=16'h3867;
aud[824]=16'h3871;
aud[825]=16'h387b;
aud[826]=16'h3886;
aud[827]=16'h3890;
aud[828]=16'h389a;
aud[829]=16'h38a4;
aud[830]=16'h38ae;
aud[831]=16'h38b8;
aud[832]=16'h38c1;
aud[833]=16'h38cb;
aud[834]=16'h38d5;
aud[835]=16'h38df;
aud[836]=16'h38e9;
aud[837]=16'h38f3;
aud[838]=16'h38fd;
aud[839]=16'h3906;
aud[840]=16'h3910;
aud[841]=16'h391a;
aud[842]=16'h3923;
aud[843]=16'h392d;
aud[844]=16'h3937;
aud[845]=16'h3940;
aud[846]=16'h394a;
aud[847]=16'h3953;
aud[848]=16'h395d;
aud[849]=16'h3966;
aud[850]=16'h3970;
aud[851]=16'h3979;
aud[852]=16'h3983;
aud[853]=16'h398c;
aud[854]=16'h3995;
aud[855]=16'h399f;
aud[856]=16'h39a8;
aud[857]=16'h39b1;
aud[858]=16'h39bb;
aud[859]=16'h39c4;
aud[860]=16'h39cd;
aud[861]=16'h39d6;
aud[862]=16'h39e0;
aud[863]=16'h39e9;
aud[864]=16'h39f2;
aud[865]=16'h39fb;
aud[866]=16'h3a04;
aud[867]=16'h3a0d;
aud[868]=16'h3a16;
aud[869]=16'h3a1f;
aud[870]=16'h3a28;
aud[871]=16'h3a31;
aud[872]=16'h3a3a;
aud[873]=16'h3a43;
aud[874]=16'h3a4c;
aud[875]=16'h3a54;
aud[876]=16'h3a5d;
aud[877]=16'h3a66;
aud[878]=16'h3a6f;
aud[879]=16'h3a78;
aud[880]=16'h3a80;
aud[881]=16'h3a89;
aud[882]=16'h3a92;
aud[883]=16'h3a9a;
aud[884]=16'h3aa3;
aud[885]=16'h3aab;
aud[886]=16'h3ab4;
aud[887]=16'h3abc;
aud[888]=16'h3ac5;
aud[889]=16'h3acd;
aud[890]=16'h3ad6;
aud[891]=16'h3ade;
aud[892]=16'h3ae7;
aud[893]=16'h3aef;
aud[894]=16'h3af7;
aud[895]=16'h3b00;
aud[896]=16'h3b08;
aud[897]=16'h3b10;
aud[898]=16'h3b19;
aud[899]=16'h3b21;
aud[900]=16'h3b29;
aud[901]=16'h3b31;
aud[902]=16'h3b39;
aud[903]=16'h3b41;
aud[904]=16'h3b4a;
aud[905]=16'h3b52;
aud[906]=16'h3b5a;
aud[907]=16'h3b62;
aud[908]=16'h3b6a;
aud[909]=16'h3b72;
aud[910]=16'h3b7a;
aud[911]=16'h3b81;
aud[912]=16'h3b89;
aud[913]=16'h3b91;
aud[914]=16'h3b99;
aud[915]=16'h3ba1;
aud[916]=16'h3ba9;
aud[917]=16'h3bb0;
aud[918]=16'h3bb8;
aud[919]=16'h3bc0;
aud[920]=16'h3bc7;
aud[921]=16'h3bcf;
aud[922]=16'h3bd7;
aud[923]=16'h3bde;
aud[924]=16'h3be6;
aud[925]=16'h3bed;
aud[926]=16'h3bf5;
aud[927]=16'h3bfc;
aud[928]=16'h3c04;
aud[929]=16'h3c0b;
aud[930]=16'h3c13;
aud[931]=16'h3c1a;
aud[932]=16'h3c21;
aud[933]=16'h3c29;
aud[934]=16'h3c30;
aud[935]=16'h3c37;
aud[936]=16'h3c3f;
aud[937]=16'h3c46;
aud[938]=16'h3c4d;
aud[939]=16'h3c54;
aud[940]=16'h3c5b;
aud[941]=16'h3c63;
aud[942]=16'h3c6a;
aud[943]=16'h3c71;
aud[944]=16'h3c78;
aud[945]=16'h3c7f;
aud[946]=16'h3c86;
aud[947]=16'h3c8d;
aud[948]=16'h3c94;
aud[949]=16'h3c9b;
aud[950]=16'h3ca1;
aud[951]=16'h3ca8;
aud[952]=16'h3caf;
aud[953]=16'h3cb6;
aud[954]=16'h3cbd;
aud[955]=16'h3cc3;
aud[956]=16'h3cca;
aud[957]=16'h3cd1;
aud[958]=16'h3cd7;
aud[959]=16'h3cde;
aud[960]=16'h3ce5;
aud[961]=16'h3ceb;
aud[962]=16'h3cf2;
aud[963]=16'h3cf8;
aud[964]=16'h3cff;
aud[965]=16'h3d05;
aud[966]=16'h3d0c;
aud[967]=16'h3d12;
aud[968]=16'h3d19;
aud[969]=16'h3d1f;
aud[970]=16'h3d25;
aud[971]=16'h3d2c;
aud[972]=16'h3d32;
aud[973]=16'h3d38;
aud[974]=16'h3d3f;
aud[975]=16'h3d45;
aud[976]=16'h3d4b;
aud[977]=16'h3d51;
aud[978]=16'h3d57;
aud[979]=16'h3d5d;
aud[980]=16'h3d63;
aud[981]=16'h3d69;
aud[982]=16'h3d6f;
aud[983]=16'h3d75;
aud[984]=16'h3d7b;
aud[985]=16'h3d81;
aud[986]=16'h3d87;
aud[987]=16'h3d8d;
aud[988]=16'h3d93;
aud[989]=16'h3d99;
aud[990]=16'h3d9f;
aud[991]=16'h3da4;
aud[992]=16'h3daa;
aud[993]=16'h3db0;
aud[994]=16'h3db6;
aud[995]=16'h3dbb;
aud[996]=16'h3dc1;
aud[997]=16'h3dc7;
aud[998]=16'h3dcc;
aud[999]=16'h3dd2;
aud[1000]=16'h3dd7;
aud[1001]=16'h3ddd;
aud[1002]=16'h3de2;
aud[1003]=16'h3de8;
aud[1004]=16'h3ded;
aud[1005]=16'h3df3;
aud[1006]=16'h3df8;
aud[1007]=16'h3dfd;
aud[1008]=16'h3e03;
aud[1009]=16'h3e08;
aud[1010]=16'h3e0d;
aud[1011]=16'h3e12;
aud[1012]=16'h3e18;
aud[1013]=16'h3e1d;
aud[1014]=16'h3e22;
aud[1015]=16'h3e27;
aud[1016]=16'h3e2c;
aud[1017]=16'h3e31;
aud[1018]=16'h3e36;
aud[1019]=16'h3e3b;
aud[1020]=16'h3e40;
aud[1021]=16'h3e45;
aud[1022]=16'h3e4a;
aud[1023]=16'h3e4f;
aud[1024]=16'h3e54;
aud[1025]=16'h3e59;
aud[1026]=16'h3e5e;
aud[1027]=16'h3e62;
aud[1028]=16'h3e67;
aud[1029]=16'h3e6c;
aud[1030]=16'h3e71;
aud[1031]=16'h3e75;
aud[1032]=16'h3e7a;
aud[1033]=16'h3e7f;
aud[1034]=16'h3e83;
aud[1035]=16'h3e88;
aud[1036]=16'h3e8c;
aud[1037]=16'h3e91;
aud[1038]=16'h3e95;
aud[1039]=16'h3e9a;
aud[1040]=16'h3e9e;
aud[1041]=16'h3ea3;
aud[1042]=16'h3ea7;
aud[1043]=16'h3eac;
aud[1044]=16'h3eb0;
aud[1045]=16'h3eb4;
aud[1046]=16'h3eb9;
aud[1047]=16'h3ebd;
aud[1048]=16'h3ec1;
aud[1049]=16'h3ec5;
aud[1050]=16'h3ec9;
aud[1051]=16'h3ecd;
aud[1052]=16'h3ed2;
aud[1053]=16'h3ed6;
aud[1054]=16'h3eda;
aud[1055]=16'h3ede;
aud[1056]=16'h3ee2;
aud[1057]=16'h3ee6;
aud[1058]=16'h3eea;
aud[1059]=16'h3eee;
aud[1060]=16'h3ef2;
aud[1061]=16'h3ef5;
aud[1062]=16'h3ef9;
aud[1063]=16'h3efd;
aud[1064]=16'h3f01;
aud[1065]=16'h3f05;
aud[1066]=16'h3f08;
aud[1067]=16'h3f0c;
aud[1068]=16'h3f10;
aud[1069]=16'h3f13;
aud[1070]=16'h3f17;
aud[1071]=16'h3f1b;
aud[1072]=16'h3f1e;
aud[1073]=16'h3f22;
aud[1074]=16'h3f25;
aud[1075]=16'h3f29;
aud[1076]=16'h3f2c;
aud[1077]=16'h3f30;
aud[1078]=16'h3f33;
aud[1079]=16'h3f36;
aud[1080]=16'h3f3a;
aud[1081]=16'h3f3d;
aud[1082]=16'h3f40;
aud[1083]=16'h3f43;
aud[1084]=16'h3f47;
aud[1085]=16'h3f4a;
aud[1086]=16'h3f4d;
aud[1087]=16'h3f50;
aud[1088]=16'h3f53;
aud[1089]=16'h3f56;
aud[1090]=16'h3f5a;
aud[1091]=16'h3f5d;
aud[1092]=16'h3f60;
aud[1093]=16'h3f63;
aud[1094]=16'h3f65;
aud[1095]=16'h3f68;
aud[1096]=16'h3f6b;
aud[1097]=16'h3f6e;
aud[1098]=16'h3f71;
aud[1099]=16'h3f74;
aud[1100]=16'h3f77;
aud[1101]=16'h3f79;
aud[1102]=16'h3f7c;
aud[1103]=16'h3f7f;
aud[1104]=16'h3f81;
aud[1105]=16'h3f84;
aud[1106]=16'h3f87;
aud[1107]=16'h3f89;
aud[1108]=16'h3f8c;
aud[1109]=16'h3f8e;
aud[1110]=16'h3f91;
aud[1111]=16'h3f93;
aud[1112]=16'h3f96;
aud[1113]=16'h3f98;
aud[1114]=16'h3f9b;
aud[1115]=16'h3f9d;
aud[1116]=16'h3f9f;
aud[1117]=16'h3fa2;
aud[1118]=16'h3fa4;
aud[1119]=16'h3fa6;
aud[1120]=16'h3fa8;
aud[1121]=16'h3fab;
aud[1122]=16'h3fad;
aud[1123]=16'h3faf;
aud[1124]=16'h3fb1;
aud[1125]=16'h3fb3;
aud[1126]=16'h3fb5;
aud[1127]=16'h3fb7;
aud[1128]=16'h3fb9;
aud[1129]=16'h3fbb;
aud[1130]=16'h3fbd;
aud[1131]=16'h3fbf;
aud[1132]=16'h3fc1;
aud[1133]=16'h3fc3;
aud[1134]=16'h3fc5;
aud[1135]=16'h3fc7;
aud[1136]=16'h3fc8;
aud[1137]=16'h3fca;
aud[1138]=16'h3fcc;
aud[1139]=16'h3fcd;
aud[1140]=16'h3fcf;
aud[1141]=16'h3fd1;
aud[1142]=16'h3fd2;
aud[1143]=16'h3fd4;
aud[1144]=16'h3fd6;
aud[1145]=16'h3fd7;
aud[1146]=16'h3fd9;
aud[1147]=16'h3fda;
aud[1148]=16'h3fdc;
aud[1149]=16'h3fdd;
aud[1150]=16'h3fde;
aud[1151]=16'h3fe0;
aud[1152]=16'h3fe1;
aud[1153]=16'h3fe2;
aud[1154]=16'h3fe4;
aud[1155]=16'h3fe5;
aud[1156]=16'h3fe6;
aud[1157]=16'h3fe7;
aud[1158]=16'h3fe8;
aud[1159]=16'h3fea;
aud[1160]=16'h3feb;
aud[1161]=16'h3fec;
aud[1162]=16'h3fed;
aud[1163]=16'h3fee;
aud[1164]=16'h3fef;
aud[1165]=16'h3ff0;
aud[1166]=16'h3ff1;
aud[1167]=16'h3ff2;
aud[1168]=16'h3ff3;
aud[1169]=16'h3ff3;
aud[1170]=16'h3ff4;
aud[1171]=16'h3ff5;
aud[1172]=16'h3ff6;
aud[1173]=16'h3ff7;
aud[1174]=16'h3ff7;
aud[1175]=16'h3ff8;
aud[1176]=16'h3ff9;
aud[1177]=16'h3ff9;
aud[1178]=16'h3ffa;
aud[1179]=16'h3ffa;
aud[1180]=16'h3ffb;
aud[1181]=16'h3ffb;
aud[1182]=16'h3ffc;
aud[1183]=16'h3ffc;
aud[1184]=16'h3ffd;
aud[1185]=16'h3ffd;
aud[1186]=16'h3ffe;
aud[1187]=16'h3ffe;
aud[1188]=16'h3ffe;
aud[1189]=16'h3fff;
aud[1190]=16'h3fff;
aud[1191]=16'h3fff;
aud[1192]=16'h3fff;
aud[1193]=16'h3fff;
aud[1194]=16'h4000;
aud[1195]=16'h4000;
aud[1196]=16'h4000;
aud[1197]=16'h4000;
aud[1198]=16'h4000;
aud[1199]=16'h4000;
aud[1200]=16'h4000;
aud[1201]=16'h4000;
aud[1202]=16'h4000;
aud[1203]=16'h4000;
aud[1204]=16'h4000;
aud[1205]=16'h3fff;
aud[1206]=16'h3fff;
aud[1207]=16'h3fff;
aud[1208]=16'h3fff;
aud[1209]=16'h3fff;
aud[1210]=16'h3ffe;
aud[1211]=16'h3ffe;
aud[1212]=16'h3ffe;
aud[1213]=16'h3ffd;
aud[1214]=16'h3ffd;
aud[1215]=16'h3ffc;
aud[1216]=16'h3ffc;
aud[1217]=16'h3ffb;
aud[1218]=16'h3ffb;
aud[1219]=16'h3ffa;
aud[1220]=16'h3ffa;
aud[1221]=16'h3ff9;
aud[1222]=16'h3ff9;
aud[1223]=16'h3ff8;
aud[1224]=16'h3ff7;
aud[1225]=16'h3ff7;
aud[1226]=16'h3ff6;
aud[1227]=16'h3ff5;
aud[1228]=16'h3ff4;
aud[1229]=16'h3ff3;
aud[1230]=16'h3ff3;
aud[1231]=16'h3ff2;
aud[1232]=16'h3ff1;
aud[1233]=16'h3ff0;
aud[1234]=16'h3fef;
aud[1235]=16'h3fee;
aud[1236]=16'h3fed;
aud[1237]=16'h3fec;
aud[1238]=16'h3feb;
aud[1239]=16'h3fea;
aud[1240]=16'h3fe8;
aud[1241]=16'h3fe7;
aud[1242]=16'h3fe6;
aud[1243]=16'h3fe5;
aud[1244]=16'h3fe4;
aud[1245]=16'h3fe2;
aud[1246]=16'h3fe1;
aud[1247]=16'h3fe0;
aud[1248]=16'h3fde;
aud[1249]=16'h3fdd;
aud[1250]=16'h3fdc;
aud[1251]=16'h3fda;
aud[1252]=16'h3fd9;
aud[1253]=16'h3fd7;
aud[1254]=16'h3fd6;
aud[1255]=16'h3fd4;
aud[1256]=16'h3fd2;
aud[1257]=16'h3fd1;
aud[1258]=16'h3fcf;
aud[1259]=16'h3fcd;
aud[1260]=16'h3fcc;
aud[1261]=16'h3fca;
aud[1262]=16'h3fc8;
aud[1263]=16'h3fc7;
aud[1264]=16'h3fc5;
aud[1265]=16'h3fc3;
aud[1266]=16'h3fc1;
aud[1267]=16'h3fbf;
aud[1268]=16'h3fbd;
aud[1269]=16'h3fbb;
aud[1270]=16'h3fb9;
aud[1271]=16'h3fb7;
aud[1272]=16'h3fb5;
aud[1273]=16'h3fb3;
aud[1274]=16'h3fb1;
aud[1275]=16'h3faf;
aud[1276]=16'h3fad;
aud[1277]=16'h3fab;
aud[1278]=16'h3fa8;
aud[1279]=16'h3fa6;
aud[1280]=16'h3fa4;
aud[1281]=16'h3fa2;
aud[1282]=16'h3f9f;
aud[1283]=16'h3f9d;
aud[1284]=16'h3f9b;
aud[1285]=16'h3f98;
aud[1286]=16'h3f96;
aud[1287]=16'h3f93;
aud[1288]=16'h3f91;
aud[1289]=16'h3f8e;
aud[1290]=16'h3f8c;
aud[1291]=16'h3f89;
aud[1292]=16'h3f87;
aud[1293]=16'h3f84;
aud[1294]=16'h3f81;
aud[1295]=16'h3f7f;
aud[1296]=16'h3f7c;
aud[1297]=16'h3f79;
aud[1298]=16'h3f77;
aud[1299]=16'h3f74;
aud[1300]=16'h3f71;
aud[1301]=16'h3f6e;
aud[1302]=16'h3f6b;
aud[1303]=16'h3f68;
aud[1304]=16'h3f65;
aud[1305]=16'h3f63;
aud[1306]=16'h3f60;
aud[1307]=16'h3f5d;
aud[1308]=16'h3f5a;
aud[1309]=16'h3f56;
aud[1310]=16'h3f53;
aud[1311]=16'h3f50;
aud[1312]=16'h3f4d;
aud[1313]=16'h3f4a;
aud[1314]=16'h3f47;
aud[1315]=16'h3f43;
aud[1316]=16'h3f40;
aud[1317]=16'h3f3d;
aud[1318]=16'h3f3a;
aud[1319]=16'h3f36;
aud[1320]=16'h3f33;
aud[1321]=16'h3f30;
aud[1322]=16'h3f2c;
aud[1323]=16'h3f29;
aud[1324]=16'h3f25;
aud[1325]=16'h3f22;
aud[1326]=16'h3f1e;
aud[1327]=16'h3f1b;
aud[1328]=16'h3f17;
aud[1329]=16'h3f13;
aud[1330]=16'h3f10;
aud[1331]=16'h3f0c;
aud[1332]=16'h3f08;
aud[1333]=16'h3f05;
aud[1334]=16'h3f01;
aud[1335]=16'h3efd;
aud[1336]=16'h3ef9;
aud[1337]=16'h3ef5;
aud[1338]=16'h3ef2;
aud[1339]=16'h3eee;
aud[1340]=16'h3eea;
aud[1341]=16'h3ee6;
aud[1342]=16'h3ee2;
aud[1343]=16'h3ede;
aud[1344]=16'h3eda;
aud[1345]=16'h3ed6;
aud[1346]=16'h3ed2;
aud[1347]=16'h3ecd;
aud[1348]=16'h3ec9;
aud[1349]=16'h3ec5;
aud[1350]=16'h3ec1;
aud[1351]=16'h3ebd;
aud[1352]=16'h3eb9;
aud[1353]=16'h3eb4;
aud[1354]=16'h3eb0;
aud[1355]=16'h3eac;
aud[1356]=16'h3ea7;
aud[1357]=16'h3ea3;
aud[1358]=16'h3e9e;
aud[1359]=16'h3e9a;
aud[1360]=16'h3e95;
aud[1361]=16'h3e91;
aud[1362]=16'h3e8c;
aud[1363]=16'h3e88;
aud[1364]=16'h3e83;
aud[1365]=16'h3e7f;
aud[1366]=16'h3e7a;
aud[1367]=16'h3e75;
aud[1368]=16'h3e71;
aud[1369]=16'h3e6c;
aud[1370]=16'h3e67;
aud[1371]=16'h3e62;
aud[1372]=16'h3e5e;
aud[1373]=16'h3e59;
aud[1374]=16'h3e54;
aud[1375]=16'h3e4f;
aud[1376]=16'h3e4a;
aud[1377]=16'h3e45;
aud[1378]=16'h3e40;
aud[1379]=16'h3e3b;
aud[1380]=16'h3e36;
aud[1381]=16'h3e31;
aud[1382]=16'h3e2c;
aud[1383]=16'h3e27;
aud[1384]=16'h3e22;
aud[1385]=16'h3e1d;
aud[1386]=16'h3e18;
aud[1387]=16'h3e12;
aud[1388]=16'h3e0d;
aud[1389]=16'h3e08;
aud[1390]=16'h3e03;
aud[1391]=16'h3dfd;
aud[1392]=16'h3df8;
aud[1393]=16'h3df3;
aud[1394]=16'h3ded;
aud[1395]=16'h3de8;
aud[1396]=16'h3de2;
aud[1397]=16'h3ddd;
aud[1398]=16'h3dd7;
aud[1399]=16'h3dd2;
aud[1400]=16'h3dcc;
aud[1401]=16'h3dc7;
aud[1402]=16'h3dc1;
aud[1403]=16'h3dbb;
aud[1404]=16'h3db6;
aud[1405]=16'h3db0;
aud[1406]=16'h3daa;
aud[1407]=16'h3da4;
aud[1408]=16'h3d9f;
aud[1409]=16'h3d99;
aud[1410]=16'h3d93;
aud[1411]=16'h3d8d;
aud[1412]=16'h3d87;
aud[1413]=16'h3d81;
aud[1414]=16'h3d7b;
aud[1415]=16'h3d75;
aud[1416]=16'h3d6f;
aud[1417]=16'h3d69;
aud[1418]=16'h3d63;
aud[1419]=16'h3d5d;
aud[1420]=16'h3d57;
aud[1421]=16'h3d51;
aud[1422]=16'h3d4b;
aud[1423]=16'h3d45;
aud[1424]=16'h3d3f;
aud[1425]=16'h3d38;
aud[1426]=16'h3d32;
aud[1427]=16'h3d2c;
aud[1428]=16'h3d25;
aud[1429]=16'h3d1f;
aud[1430]=16'h3d19;
aud[1431]=16'h3d12;
aud[1432]=16'h3d0c;
aud[1433]=16'h3d05;
aud[1434]=16'h3cff;
aud[1435]=16'h3cf8;
aud[1436]=16'h3cf2;
aud[1437]=16'h3ceb;
aud[1438]=16'h3ce5;
aud[1439]=16'h3cde;
aud[1440]=16'h3cd7;
aud[1441]=16'h3cd1;
aud[1442]=16'h3cca;
aud[1443]=16'h3cc3;
aud[1444]=16'h3cbd;
aud[1445]=16'h3cb6;
aud[1446]=16'h3caf;
aud[1447]=16'h3ca8;
aud[1448]=16'h3ca1;
aud[1449]=16'h3c9b;
aud[1450]=16'h3c94;
aud[1451]=16'h3c8d;
aud[1452]=16'h3c86;
aud[1453]=16'h3c7f;
aud[1454]=16'h3c78;
aud[1455]=16'h3c71;
aud[1456]=16'h3c6a;
aud[1457]=16'h3c63;
aud[1458]=16'h3c5b;
aud[1459]=16'h3c54;
aud[1460]=16'h3c4d;
aud[1461]=16'h3c46;
aud[1462]=16'h3c3f;
aud[1463]=16'h3c37;
aud[1464]=16'h3c30;
aud[1465]=16'h3c29;
aud[1466]=16'h3c21;
aud[1467]=16'h3c1a;
aud[1468]=16'h3c13;
aud[1469]=16'h3c0b;
aud[1470]=16'h3c04;
aud[1471]=16'h3bfc;
aud[1472]=16'h3bf5;
aud[1473]=16'h3bed;
aud[1474]=16'h3be6;
aud[1475]=16'h3bde;
aud[1476]=16'h3bd7;
aud[1477]=16'h3bcf;
aud[1478]=16'h3bc7;
aud[1479]=16'h3bc0;
aud[1480]=16'h3bb8;
aud[1481]=16'h3bb0;
aud[1482]=16'h3ba9;
aud[1483]=16'h3ba1;
aud[1484]=16'h3b99;
aud[1485]=16'h3b91;
aud[1486]=16'h3b89;
aud[1487]=16'h3b81;
aud[1488]=16'h3b7a;
aud[1489]=16'h3b72;
aud[1490]=16'h3b6a;
aud[1491]=16'h3b62;
aud[1492]=16'h3b5a;
aud[1493]=16'h3b52;
aud[1494]=16'h3b4a;
aud[1495]=16'h3b41;
aud[1496]=16'h3b39;
aud[1497]=16'h3b31;
aud[1498]=16'h3b29;
aud[1499]=16'h3b21;
aud[1500]=16'h3b19;
aud[1501]=16'h3b10;
aud[1502]=16'h3b08;
aud[1503]=16'h3b00;
aud[1504]=16'h3af7;
aud[1505]=16'h3aef;
aud[1506]=16'h3ae7;
aud[1507]=16'h3ade;
aud[1508]=16'h3ad6;
aud[1509]=16'h3acd;
aud[1510]=16'h3ac5;
aud[1511]=16'h3abc;
aud[1512]=16'h3ab4;
aud[1513]=16'h3aab;
aud[1514]=16'h3aa3;
aud[1515]=16'h3a9a;
aud[1516]=16'h3a92;
aud[1517]=16'h3a89;
aud[1518]=16'h3a80;
aud[1519]=16'h3a78;
aud[1520]=16'h3a6f;
aud[1521]=16'h3a66;
aud[1522]=16'h3a5d;
aud[1523]=16'h3a54;
aud[1524]=16'h3a4c;
aud[1525]=16'h3a43;
aud[1526]=16'h3a3a;
aud[1527]=16'h3a31;
aud[1528]=16'h3a28;
aud[1529]=16'h3a1f;
aud[1530]=16'h3a16;
aud[1531]=16'h3a0d;
aud[1532]=16'h3a04;
aud[1533]=16'h39fb;
aud[1534]=16'h39f2;
aud[1535]=16'h39e9;
aud[1536]=16'h39e0;
aud[1537]=16'h39d6;
aud[1538]=16'h39cd;
aud[1539]=16'h39c4;
aud[1540]=16'h39bb;
aud[1541]=16'h39b1;
aud[1542]=16'h39a8;
aud[1543]=16'h399f;
aud[1544]=16'h3995;
aud[1545]=16'h398c;
aud[1546]=16'h3983;
aud[1547]=16'h3979;
aud[1548]=16'h3970;
aud[1549]=16'h3966;
aud[1550]=16'h395d;
aud[1551]=16'h3953;
aud[1552]=16'h394a;
aud[1553]=16'h3940;
aud[1554]=16'h3937;
aud[1555]=16'h392d;
aud[1556]=16'h3923;
aud[1557]=16'h391a;
aud[1558]=16'h3910;
aud[1559]=16'h3906;
aud[1560]=16'h38fd;
aud[1561]=16'h38f3;
aud[1562]=16'h38e9;
aud[1563]=16'h38df;
aud[1564]=16'h38d5;
aud[1565]=16'h38cb;
aud[1566]=16'h38c1;
aud[1567]=16'h38b8;
aud[1568]=16'h38ae;
aud[1569]=16'h38a4;
aud[1570]=16'h389a;
aud[1571]=16'h3890;
aud[1572]=16'h3886;
aud[1573]=16'h387b;
aud[1574]=16'h3871;
aud[1575]=16'h3867;
aud[1576]=16'h385d;
aud[1577]=16'h3853;
aud[1578]=16'h3849;
aud[1579]=16'h383f;
aud[1580]=16'h3834;
aud[1581]=16'h382a;
aud[1582]=16'h3820;
aud[1583]=16'h3815;
aud[1584]=16'h380b;
aud[1585]=16'h3801;
aud[1586]=16'h37f6;
aud[1587]=16'h37ec;
aud[1588]=16'h37e1;
aud[1589]=16'h37d7;
aud[1590]=16'h37cc;
aud[1591]=16'h37c2;
aud[1592]=16'h37b7;
aud[1593]=16'h37ad;
aud[1594]=16'h37a2;
aud[1595]=16'h3798;
aud[1596]=16'h378d;
aud[1597]=16'h3782;
aud[1598]=16'h3778;
aud[1599]=16'h376d;
aud[1600]=16'h3762;
aud[1601]=16'h3757;
aud[1602]=16'h374d;
aud[1603]=16'h3742;
aud[1604]=16'h3737;
aud[1605]=16'h372c;
aud[1606]=16'h3721;
aud[1607]=16'h3716;
aud[1608]=16'h370b;
aud[1609]=16'h3701;
aud[1610]=16'h36f6;
aud[1611]=16'h36eb;
aud[1612]=16'h36e0;
aud[1613]=16'h36d4;
aud[1614]=16'h36c9;
aud[1615]=16'h36be;
aud[1616]=16'h36b3;
aud[1617]=16'h36a8;
aud[1618]=16'h369d;
aud[1619]=16'h3692;
aud[1620]=16'h3686;
aud[1621]=16'h367b;
aud[1622]=16'h3670;
aud[1623]=16'h3665;
aud[1624]=16'h3659;
aud[1625]=16'h364e;
aud[1626]=16'h3643;
aud[1627]=16'h3637;
aud[1628]=16'h362c;
aud[1629]=16'h3620;
aud[1630]=16'h3615;
aud[1631]=16'h3609;
aud[1632]=16'h35fe;
aud[1633]=16'h35f2;
aud[1634]=16'h35e7;
aud[1635]=16'h35db;
aud[1636]=16'h35d0;
aud[1637]=16'h35c4;
aud[1638]=16'h35b8;
aud[1639]=16'h35ad;
aud[1640]=16'h35a1;
aud[1641]=16'h3595;
aud[1642]=16'h358a;
aud[1643]=16'h357e;
aud[1644]=16'h3572;
aud[1645]=16'h3566;
aud[1646]=16'h355a;
aud[1647]=16'h354f;
aud[1648]=16'h3543;
aud[1649]=16'h3537;
aud[1650]=16'h352b;
aud[1651]=16'h351f;
aud[1652]=16'h3513;
aud[1653]=16'h3507;
aud[1654]=16'h34fb;
aud[1655]=16'h34ef;
aud[1656]=16'h34e3;
aud[1657]=16'h34d7;
aud[1658]=16'h34cb;
aud[1659]=16'h34be;
aud[1660]=16'h34b2;
aud[1661]=16'h34a6;
aud[1662]=16'h349a;
aud[1663]=16'h348e;
aud[1664]=16'h3481;
aud[1665]=16'h3475;
aud[1666]=16'h3469;
aud[1667]=16'h345d;
aud[1668]=16'h3450;
aud[1669]=16'h3444;
aud[1670]=16'h3437;
aud[1671]=16'h342b;
aud[1672]=16'h341f;
aud[1673]=16'h3412;
aud[1674]=16'h3406;
aud[1675]=16'h33f9;
aud[1676]=16'h33ed;
aud[1677]=16'h33e0;
aud[1678]=16'h33d4;
aud[1679]=16'h33c7;
aud[1680]=16'h33ba;
aud[1681]=16'h33ae;
aud[1682]=16'h33a1;
aud[1683]=16'h3394;
aud[1684]=16'h3388;
aud[1685]=16'h337b;
aud[1686]=16'h336e;
aud[1687]=16'h3361;
aud[1688]=16'h3355;
aud[1689]=16'h3348;
aud[1690]=16'h333b;
aud[1691]=16'h332e;
aud[1692]=16'h3321;
aud[1693]=16'h3314;
aud[1694]=16'h3307;
aud[1695]=16'h32fa;
aud[1696]=16'h32ed;
aud[1697]=16'h32e0;
aud[1698]=16'h32d3;
aud[1699]=16'h32c6;
aud[1700]=16'h32b9;
aud[1701]=16'h32ac;
aud[1702]=16'h329f;
aud[1703]=16'h3292;
aud[1704]=16'h3285;
aud[1705]=16'h3278;
aud[1706]=16'h326a;
aud[1707]=16'h325d;
aud[1708]=16'h3250;
aud[1709]=16'h3243;
aud[1710]=16'h3235;
aud[1711]=16'h3228;
aud[1712]=16'h321b;
aud[1713]=16'h320d;
aud[1714]=16'h3200;
aud[1715]=16'h31f3;
aud[1716]=16'h31e5;
aud[1717]=16'h31d8;
aud[1718]=16'h31ca;
aud[1719]=16'h31bd;
aud[1720]=16'h31af;
aud[1721]=16'h31a2;
aud[1722]=16'h3194;
aud[1723]=16'h3187;
aud[1724]=16'h3179;
aud[1725]=16'h316b;
aud[1726]=16'h315e;
aud[1727]=16'h3150;
aud[1728]=16'h3142;
aud[1729]=16'h3135;
aud[1730]=16'h3127;
aud[1731]=16'h3119;
aud[1732]=16'h310b;
aud[1733]=16'h30fe;
aud[1734]=16'h30f0;
aud[1735]=16'h30e2;
aud[1736]=16'h30d4;
aud[1737]=16'h30c6;
aud[1738]=16'h30b8;
aud[1739]=16'h30aa;
aud[1740]=16'h309d;
aud[1741]=16'h308f;
aud[1742]=16'h3081;
aud[1743]=16'h3073;
aud[1744]=16'h3065;
aud[1745]=16'h3057;
aud[1746]=16'h3048;
aud[1747]=16'h303a;
aud[1748]=16'h302c;
aud[1749]=16'h301e;
aud[1750]=16'h3010;
aud[1751]=16'h3002;
aud[1752]=16'h2ff4;
aud[1753]=16'h2fe5;
aud[1754]=16'h2fd7;
aud[1755]=16'h2fc9;
aud[1756]=16'h2fbb;
aud[1757]=16'h2fac;
aud[1758]=16'h2f9e;
aud[1759]=16'h2f90;
aud[1760]=16'h2f81;
aud[1761]=16'h2f73;
aud[1762]=16'h2f65;
aud[1763]=16'h2f56;
aud[1764]=16'h2f48;
aud[1765]=16'h2f39;
aud[1766]=16'h2f2b;
aud[1767]=16'h2f1c;
aud[1768]=16'h2f0e;
aud[1769]=16'h2eff;
aud[1770]=16'h2ef1;
aud[1771]=16'h2ee2;
aud[1772]=16'h2ed3;
aud[1773]=16'h2ec5;
aud[1774]=16'h2eb6;
aud[1775]=16'h2ea7;
aud[1776]=16'h2e99;
aud[1777]=16'h2e8a;
aud[1778]=16'h2e7b;
aud[1779]=16'h2e6d;
aud[1780]=16'h2e5e;
aud[1781]=16'h2e4f;
aud[1782]=16'h2e40;
aud[1783]=16'h2e31;
aud[1784]=16'h2e22;
aud[1785]=16'h2e14;
aud[1786]=16'h2e05;
aud[1787]=16'h2df6;
aud[1788]=16'h2de7;
aud[1789]=16'h2dd8;
aud[1790]=16'h2dc9;
aud[1791]=16'h2dba;
aud[1792]=16'h2dab;
aud[1793]=16'h2d9c;
aud[1794]=16'h2d8d;
aud[1795]=16'h2d7e;
aud[1796]=16'h2d6f;
aud[1797]=16'h2d60;
aud[1798]=16'h2d50;
aud[1799]=16'h2d41;
aud[1800]=16'h2d32;
aud[1801]=16'h2d23;
aud[1802]=16'h2d14;
aud[1803]=16'h2d04;
aud[1804]=16'h2cf5;
aud[1805]=16'h2ce6;
aud[1806]=16'h2cd7;
aud[1807]=16'h2cc7;
aud[1808]=16'h2cb8;
aud[1809]=16'h2ca9;
aud[1810]=16'h2c99;
aud[1811]=16'h2c8a;
aud[1812]=16'h2c7a;
aud[1813]=16'h2c6b;
aud[1814]=16'h2c5c;
aud[1815]=16'h2c4c;
aud[1816]=16'h2c3d;
aud[1817]=16'h2c2d;
aud[1818]=16'h2c1e;
aud[1819]=16'h2c0e;
aud[1820]=16'h2bfe;
aud[1821]=16'h2bef;
aud[1822]=16'h2bdf;
aud[1823]=16'h2bd0;
aud[1824]=16'h2bc0;
aud[1825]=16'h2bb0;
aud[1826]=16'h2ba1;
aud[1827]=16'h2b91;
aud[1828]=16'h2b81;
aud[1829]=16'h2b71;
aud[1830]=16'h2b62;
aud[1831]=16'h2b52;
aud[1832]=16'h2b42;
aud[1833]=16'h2b32;
aud[1834]=16'h2b22;
aud[1835]=16'h2b13;
aud[1836]=16'h2b03;
aud[1837]=16'h2af3;
aud[1838]=16'h2ae3;
aud[1839]=16'h2ad3;
aud[1840]=16'h2ac3;
aud[1841]=16'h2ab3;
aud[1842]=16'h2aa3;
aud[1843]=16'h2a93;
aud[1844]=16'h2a83;
aud[1845]=16'h2a73;
aud[1846]=16'h2a63;
aud[1847]=16'h2a53;
aud[1848]=16'h2a43;
aud[1849]=16'h2a33;
aud[1850]=16'h2a23;
aud[1851]=16'h2a12;
aud[1852]=16'h2a02;
aud[1853]=16'h29f2;
aud[1854]=16'h29e2;
aud[1855]=16'h29d2;
aud[1856]=16'h29c1;
aud[1857]=16'h29b1;
aud[1858]=16'h29a1;
aud[1859]=16'h2991;
aud[1860]=16'h2980;
aud[1861]=16'h2970;
aud[1862]=16'h2960;
aud[1863]=16'h294f;
aud[1864]=16'h293f;
aud[1865]=16'h292e;
aud[1866]=16'h291e;
aud[1867]=16'h290e;
aud[1868]=16'h28fd;
aud[1869]=16'h28ed;
aud[1870]=16'h28dc;
aud[1871]=16'h28cc;
aud[1872]=16'h28bb;
aud[1873]=16'h28aa;
aud[1874]=16'h289a;
aud[1875]=16'h2889;
aud[1876]=16'h2879;
aud[1877]=16'h2868;
aud[1878]=16'h2857;
aud[1879]=16'h2847;
aud[1880]=16'h2836;
aud[1881]=16'h2825;
aud[1882]=16'h2815;
aud[1883]=16'h2804;
aud[1884]=16'h27f3;
aud[1885]=16'h27e2;
aud[1886]=16'h27d2;
aud[1887]=16'h27c1;
aud[1888]=16'h27b0;
aud[1889]=16'h279f;
aud[1890]=16'h278e;
aud[1891]=16'h277e;
aud[1892]=16'h276d;
aud[1893]=16'h275c;
aud[1894]=16'h274b;
aud[1895]=16'h273a;
aud[1896]=16'h2729;
aud[1897]=16'h2718;
aud[1898]=16'h2707;
aud[1899]=16'h26f6;
aud[1900]=16'h26e5;
aud[1901]=16'h26d4;
aud[1902]=16'h26c3;
aud[1903]=16'h26b2;
aud[1904]=16'h26a1;
aud[1905]=16'h2690;
aud[1906]=16'h267e;
aud[1907]=16'h266d;
aud[1908]=16'h265c;
aud[1909]=16'h264b;
aud[1910]=16'h263a;
aud[1911]=16'h2629;
aud[1912]=16'h2617;
aud[1913]=16'h2606;
aud[1914]=16'h25f5;
aud[1915]=16'h25e4;
aud[1916]=16'h25d2;
aud[1917]=16'h25c1;
aud[1918]=16'h25b0;
aud[1919]=16'h259e;
aud[1920]=16'h258d;
aud[1921]=16'h257c;
aud[1922]=16'h256a;
aud[1923]=16'h2559;
aud[1924]=16'h2547;
aud[1925]=16'h2536;
aud[1926]=16'h2524;
aud[1927]=16'h2513;
aud[1928]=16'h2501;
aud[1929]=16'h24f0;
aud[1930]=16'h24de;
aud[1931]=16'h24cd;
aud[1932]=16'h24bb;
aud[1933]=16'h24aa;
aud[1934]=16'h2498;
aud[1935]=16'h2487;
aud[1936]=16'h2475;
aud[1937]=16'h2463;
aud[1938]=16'h2452;
aud[1939]=16'h2440;
aud[1940]=16'h242e;
aud[1941]=16'h241d;
aud[1942]=16'h240b;
aud[1943]=16'h23f9;
aud[1944]=16'h23e7;
aud[1945]=16'h23d6;
aud[1946]=16'h23c4;
aud[1947]=16'h23b2;
aud[1948]=16'h23a0;
aud[1949]=16'h238e;
aud[1950]=16'h237d;
aud[1951]=16'h236b;
aud[1952]=16'h2359;
aud[1953]=16'h2347;
aud[1954]=16'h2335;
aud[1955]=16'h2323;
aud[1956]=16'h2311;
aud[1957]=16'h22ff;
aud[1958]=16'h22ed;
aud[1959]=16'h22db;
aud[1960]=16'h22c9;
aud[1961]=16'h22b7;
aud[1962]=16'h22a5;
aud[1963]=16'h2293;
aud[1964]=16'h2281;
aud[1965]=16'h226f;
aud[1966]=16'h225d;
aud[1967]=16'h224b;
aud[1968]=16'h2239;
aud[1969]=16'h2227;
aud[1970]=16'h2215;
aud[1971]=16'h2202;
aud[1972]=16'h21f0;
aud[1973]=16'h21de;
aud[1974]=16'h21cc;
aud[1975]=16'h21ba;
aud[1976]=16'h21a7;
aud[1977]=16'h2195;
aud[1978]=16'h2183;
aud[1979]=16'h2171;
aud[1980]=16'h215e;
aud[1981]=16'h214c;
aud[1982]=16'h213a;
aud[1983]=16'h2127;
aud[1984]=16'h2115;
aud[1985]=16'h2103;
aud[1986]=16'h20f0;
aud[1987]=16'h20de;
aud[1988]=16'h20cb;
aud[1989]=16'h20b9;
aud[1990]=16'h20a7;
aud[1991]=16'h2094;
aud[1992]=16'h2082;
aud[1993]=16'h206f;
aud[1994]=16'h205d;
aud[1995]=16'h204a;
aud[1996]=16'h2038;
aud[1997]=16'h2025;
aud[1998]=16'h2013;
aud[1999]=16'h2000;
aud[2000]=16'h1fed;
aud[2001]=16'h1fdb;
aud[2002]=16'h1fc8;
aud[2003]=16'h1fb6;
aud[2004]=16'h1fa3;
aud[2005]=16'h1f90;
aud[2006]=16'h1f7e;
aud[2007]=16'h1f6b;
aud[2008]=16'h1f58;
aud[2009]=16'h1f46;
aud[2010]=16'h1f33;
aud[2011]=16'h1f20;
aud[2012]=16'h1f0d;
aud[2013]=16'h1efb;
aud[2014]=16'h1ee8;
aud[2015]=16'h1ed5;
aud[2016]=16'h1ec2;
aud[2017]=16'h1eaf;
aud[2018]=16'h1e9d;
aud[2019]=16'h1e8a;
aud[2020]=16'h1e77;
aud[2021]=16'h1e64;
aud[2022]=16'h1e51;
aud[2023]=16'h1e3e;
aud[2024]=16'h1e2b;
aud[2025]=16'h1e18;
aud[2026]=16'h1e06;
aud[2027]=16'h1df3;
aud[2028]=16'h1de0;
aud[2029]=16'h1dcd;
aud[2030]=16'h1dba;
aud[2031]=16'h1da7;
aud[2032]=16'h1d94;
aud[2033]=16'h1d81;
aud[2034]=16'h1d6e;
aud[2035]=16'h1d5b;
aud[2036]=16'h1d47;
aud[2037]=16'h1d34;
aud[2038]=16'h1d21;
aud[2039]=16'h1d0e;
aud[2040]=16'h1cfb;
aud[2041]=16'h1ce8;
aud[2042]=16'h1cd5;
aud[2043]=16'h1cc2;
aud[2044]=16'h1cae;
aud[2045]=16'h1c9b;
aud[2046]=16'h1c88;
aud[2047]=16'h1c75;
aud[2048]=16'h1c62;
aud[2049]=16'h1c4e;
aud[2050]=16'h1c3b;
aud[2051]=16'h1c28;
aud[2052]=16'h1c15;
aud[2053]=16'h1c01;
aud[2054]=16'h1bee;
aud[2055]=16'h1bdb;
aud[2056]=16'h1bc8;
aud[2057]=16'h1bb4;
aud[2058]=16'h1ba1;
aud[2059]=16'h1b8d;
aud[2060]=16'h1b7a;
aud[2061]=16'h1b67;
aud[2062]=16'h1b53;
aud[2063]=16'h1b40;
aud[2064]=16'h1b2d;
aud[2065]=16'h1b19;
aud[2066]=16'h1b06;
aud[2067]=16'h1af2;
aud[2068]=16'h1adf;
aud[2069]=16'h1acb;
aud[2070]=16'h1ab8;
aud[2071]=16'h1aa4;
aud[2072]=16'h1a91;
aud[2073]=16'h1a7d;
aud[2074]=16'h1a6a;
aud[2075]=16'h1a56;
aud[2076]=16'h1a43;
aud[2077]=16'h1a2f;
aud[2078]=16'h1a1c;
aud[2079]=16'h1a08;
aud[2080]=16'h19f4;
aud[2081]=16'h19e1;
aud[2082]=16'h19cd;
aud[2083]=16'h19ba;
aud[2084]=16'h19a6;
aud[2085]=16'h1992;
aud[2086]=16'h197f;
aud[2087]=16'h196b;
aud[2088]=16'h1957;
aud[2089]=16'h1943;
aud[2090]=16'h1930;
aud[2091]=16'h191c;
aud[2092]=16'h1908;
aud[2093]=16'h18f5;
aud[2094]=16'h18e1;
aud[2095]=16'h18cd;
aud[2096]=16'h18b9;
aud[2097]=16'h18a5;
aud[2098]=16'h1892;
aud[2099]=16'h187e;
aud[2100]=16'h186a;
aud[2101]=16'h1856;
aud[2102]=16'h1842;
aud[2103]=16'h182f;
aud[2104]=16'h181b;
aud[2105]=16'h1807;
aud[2106]=16'h17f3;
aud[2107]=16'h17df;
aud[2108]=16'h17cb;
aud[2109]=16'h17b7;
aud[2110]=16'h17a3;
aud[2111]=16'h178f;
aud[2112]=16'h177b;
aud[2113]=16'h1767;
aud[2114]=16'h1753;
aud[2115]=16'h1740;
aud[2116]=16'h172c;
aud[2117]=16'h1718;
aud[2118]=16'h1704;
aud[2119]=16'h16f0;
aud[2120]=16'h16db;
aud[2121]=16'h16c7;
aud[2122]=16'h16b3;
aud[2123]=16'h169f;
aud[2124]=16'h168b;
aud[2125]=16'h1677;
aud[2126]=16'h1663;
aud[2127]=16'h164f;
aud[2128]=16'h163b;
aud[2129]=16'h1627;
aud[2130]=16'h1613;
aud[2131]=16'h15ff;
aud[2132]=16'h15ea;
aud[2133]=16'h15d6;
aud[2134]=16'h15c2;
aud[2135]=16'h15ae;
aud[2136]=16'h159a;
aud[2137]=16'h1586;
aud[2138]=16'h1571;
aud[2139]=16'h155d;
aud[2140]=16'h1549;
aud[2141]=16'h1535;
aud[2142]=16'h1520;
aud[2143]=16'h150c;
aud[2144]=16'h14f8;
aud[2145]=16'h14e4;
aud[2146]=16'h14cf;
aud[2147]=16'h14bb;
aud[2148]=16'h14a7;
aud[2149]=16'h1492;
aud[2150]=16'h147e;
aud[2151]=16'h146a;
aud[2152]=16'h1455;
aud[2153]=16'h1441;
aud[2154]=16'h142d;
aud[2155]=16'h1418;
aud[2156]=16'h1404;
aud[2157]=16'h13f0;
aud[2158]=16'h13db;
aud[2159]=16'h13c7;
aud[2160]=16'h13b3;
aud[2161]=16'h139e;
aud[2162]=16'h138a;
aud[2163]=16'h1375;
aud[2164]=16'h1361;
aud[2165]=16'h134c;
aud[2166]=16'h1338;
aud[2167]=16'h1323;
aud[2168]=16'h130f;
aud[2169]=16'h12fb;
aud[2170]=16'h12e6;
aud[2171]=16'h12d2;
aud[2172]=16'h12bd;
aud[2173]=16'h12a9;
aud[2174]=16'h1294;
aud[2175]=16'h127f;
aud[2176]=16'h126b;
aud[2177]=16'h1256;
aud[2178]=16'h1242;
aud[2179]=16'h122d;
aud[2180]=16'h1219;
aud[2181]=16'h1204;
aud[2182]=16'h11f0;
aud[2183]=16'h11db;
aud[2184]=16'h11c6;
aud[2185]=16'h11b2;
aud[2186]=16'h119d;
aud[2187]=16'h1189;
aud[2188]=16'h1174;
aud[2189]=16'h115f;
aud[2190]=16'h114b;
aud[2191]=16'h1136;
aud[2192]=16'h1121;
aud[2193]=16'h110d;
aud[2194]=16'h10f8;
aud[2195]=16'h10e3;
aud[2196]=16'h10cf;
aud[2197]=16'h10ba;
aud[2198]=16'h10a5;
aud[2199]=16'h1090;
aud[2200]=16'h107c;
aud[2201]=16'h1067;
aud[2202]=16'h1052;
aud[2203]=16'h103e;
aud[2204]=16'h1029;
aud[2205]=16'h1014;
aud[2206]=16'hfff;
aud[2207]=16'hfeb;
aud[2208]=16'hfd6;
aud[2209]=16'hfc1;
aud[2210]=16'hfac;
aud[2211]=16'hf97;
aud[2212]=16'hf83;
aud[2213]=16'hf6e;
aud[2214]=16'hf59;
aud[2215]=16'hf44;
aud[2216]=16'hf2f;
aud[2217]=16'hf1a;
aud[2218]=16'hf06;
aud[2219]=16'hef1;
aud[2220]=16'hedc;
aud[2221]=16'hec7;
aud[2222]=16'heb2;
aud[2223]=16'he9d;
aud[2224]=16'he88;
aud[2225]=16'he74;
aud[2226]=16'he5f;
aud[2227]=16'he4a;
aud[2228]=16'he35;
aud[2229]=16'he20;
aud[2230]=16'he0b;
aud[2231]=16'hdf6;
aud[2232]=16'hde1;
aud[2233]=16'hdcc;
aud[2234]=16'hdb7;
aud[2235]=16'hda2;
aud[2236]=16'hd8d;
aud[2237]=16'hd78;
aud[2238]=16'hd63;
aud[2239]=16'hd4e;
aud[2240]=16'hd39;
aud[2241]=16'hd24;
aud[2242]=16'hd0f;
aud[2243]=16'hcfa;
aud[2244]=16'hce5;
aud[2245]=16'hcd0;
aud[2246]=16'hcbb;
aud[2247]=16'hca6;
aud[2248]=16'hc91;
aud[2249]=16'hc7c;
aud[2250]=16'hc67;
aud[2251]=16'hc52;
aud[2252]=16'hc3d;
aud[2253]=16'hc28;
aud[2254]=16'hc13;
aud[2255]=16'hbfe;
aud[2256]=16'hbe9;
aud[2257]=16'hbd4;
aud[2258]=16'hbbf;
aud[2259]=16'hbaa;
aud[2260]=16'hb95;
aud[2261]=16'hb80;
aud[2262]=16'hb6a;
aud[2263]=16'hb55;
aud[2264]=16'hb40;
aud[2265]=16'hb2b;
aud[2266]=16'hb16;
aud[2267]=16'hb01;
aud[2268]=16'haec;
aud[2269]=16'had7;
aud[2270]=16'hac1;
aud[2271]=16'haac;
aud[2272]=16'ha97;
aud[2273]=16'ha82;
aud[2274]=16'ha6d;
aud[2275]=16'ha58;
aud[2276]=16'ha43;
aud[2277]=16'ha2d;
aud[2278]=16'ha18;
aud[2279]=16'ha03;
aud[2280]=16'h9ee;
aud[2281]=16'h9d9;
aud[2282]=16'h9c3;
aud[2283]=16'h9ae;
aud[2284]=16'h999;
aud[2285]=16'h984;
aud[2286]=16'h96f;
aud[2287]=16'h959;
aud[2288]=16'h944;
aud[2289]=16'h92f;
aud[2290]=16'h91a;
aud[2291]=16'h905;
aud[2292]=16'h8ef;
aud[2293]=16'h8da;
aud[2294]=16'h8c5;
aud[2295]=16'h8b0;
aud[2296]=16'h89a;
aud[2297]=16'h885;
aud[2298]=16'h870;
aud[2299]=16'h85b;
aud[2300]=16'h845;
aud[2301]=16'h830;
aud[2302]=16'h81b;
aud[2303]=16'h805;
aud[2304]=16'h7f0;
aud[2305]=16'h7db;
aud[2306]=16'h7c6;
aud[2307]=16'h7b0;
aud[2308]=16'h79b;
aud[2309]=16'h786;
aud[2310]=16'h770;
aud[2311]=16'h75b;
aud[2312]=16'h746;
aud[2313]=16'h731;
aud[2314]=16'h71b;
aud[2315]=16'h706;
aud[2316]=16'h6f1;
aud[2317]=16'h6db;
aud[2318]=16'h6c6;
aud[2319]=16'h6b1;
aud[2320]=16'h69b;
aud[2321]=16'h686;
aud[2322]=16'h671;
aud[2323]=16'h65b;
aud[2324]=16'h646;
aud[2325]=16'h631;
aud[2326]=16'h61b;
aud[2327]=16'h606;
aud[2328]=16'h5f1;
aud[2329]=16'h5db;
aud[2330]=16'h5c6;
aud[2331]=16'h5b0;
aud[2332]=16'h59b;
aud[2333]=16'h586;
aud[2334]=16'h570;
aud[2335]=16'h55b;
aud[2336]=16'h546;
aud[2337]=16'h530;
aud[2338]=16'h51b;
aud[2339]=16'h505;
aud[2340]=16'h4f0;
aud[2341]=16'h4db;
aud[2342]=16'h4c5;
aud[2343]=16'h4b0;
aud[2344]=16'h49b;
aud[2345]=16'h485;
aud[2346]=16'h470;
aud[2347]=16'h45a;
aud[2348]=16'h445;
aud[2349]=16'h430;
aud[2350]=16'h41a;
aud[2351]=16'h405;
aud[2352]=16'h3ef;
aud[2353]=16'h3da;
aud[2354]=16'h3c5;
aud[2355]=16'h3af;
aud[2356]=16'h39a;
aud[2357]=16'h384;
aud[2358]=16'h36f;
aud[2359]=16'h359;
aud[2360]=16'h344;
aud[2361]=16'h32f;
aud[2362]=16'h319;
aud[2363]=16'h304;
aud[2364]=16'h2ee;
aud[2365]=16'h2d9;
aud[2366]=16'h2c4;
aud[2367]=16'h2ae;
aud[2368]=16'h299;
aud[2369]=16'h283;
aud[2370]=16'h26e;
aud[2371]=16'h258;
aud[2372]=16'h243;
aud[2373]=16'h22e;
aud[2374]=16'h218;
aud[2375]=16'h203;
aud[2376]=16'h1ed;
aud[2377]=16'h1d8;
aud[2378]=16'h1c2;
aud[2379]=16'h1ad;
aud[2380]=16'h197;
aud[2381]=16'h182;
aud[2382]=16'h16d;
aud[2383]=16'h157;
aud[2384]=16'h142;
aud[2385]=16'h12c;
aud[2386]=16'h117;
aud[2387]=16'h101;
aud[2388]=16'hec;
aud[2389]=16'hd6;
aud[2390]=16'hc1;
aud[2391]=16'hac;
aud[2392]=16'h96;
aud[2393]=16'h81;
aud[2394]=16'h6b;
aud[2395]=16'h56;
aud[2396]=16'h40;
aud[2397]=16'h2b;
aud[2398]=16'h15;
aud[2399]=16'h0;
aud[2400]=16'hffeb;
aud[2401]=16'hffd5;
aud[2402]=16'hffc0;
aud[2403]=16'hffaa;
aud[2404]=16'hff95;
aud[2405]=16'hff7f;
aud[2406]=16'hff6a;
aud[2407]=16'hff54;
aud[2408]=16'hff3f;
aud[2409]=16'hff2a;
aud[2410]=16'hff14;
aud[2411]=16'hfeff;
aud[2412]=16'hfee9;
aud[2413]=16'hfed4;
aud[2414]=16'hfebe;
aud[2415]=16'hfea9;
aud[2416]=16'hfe93;
aud[2417]=16'hfe7e;
aud[2418]=16'hfe69;
aud[2419]=16'hfe53;
aud[2420]=16'hfe3e;
aud[2421]=16'hfe28;
aud[2422]=16'hfe13;
aud[2423]=16'hfdfd;
aud[2424]=16'hfde8;
aud[2425]=16'hfdd2;
aud[2426]=16'hfdbd;
aud[2427]=16'hfda8;
aud[2428]=16'hfd92;
aud[2429]=16'hfd7d;
aud[2430]=16'hfd67;
aud[2431]=16'hfd52;
aud[2432]=16'hfd3c;
aud[2433]=16'hfd27;
aud[2434]=16'hfd12;
aud[2435]=16'hfcfc;
aud[2436]=16'hfce7;
aud[2437]=16'hfcd1;
aud[2438]=16'hfcbc;
aud[2439]=16'hfca7;
aud[2440]=16'hfc91;
aud[2441]=16'hfc7c;
aud[2442]=16'hfc66;
aud[2443]=16'hfc51;
aud[2444]=16'hfc3b;
aud[2445]=16'hfc26;
aud[2446]=16'hfc11;
aud[2447]=16'hfbfb;
aud[2448]=16'hfbe6;
aud[2449]=16'hfbd0;
aud[2450]=16'hfbbb;
aud[2451]=16'hfba6;
aud[2452]=16'hfb90;
aud[2453]=16'hfb7b;
aud[2454]=16'hfb65;
aud[2455]=16'hfb50;
aud[2456]=16'hfb3b;
aud[2457]=16'hfb25;
aud[2458]=16'hfb10;
aud[2459]=16'hfafb;
aud[2460]=16'hfae5;
aud[2461]=16'hfad0;
aud[2462]=16'hfaba;
aud[2463]=16'hfaa5;
aud[2464]=16'hfa90;
aud[2465]=16'hfa7a;
aud[2466]=16'hfa65;
aud[2467]=16'hfa50;
aud[2468]=16'hfa3a;
aud[2469]=16'hfa25;
aud[2470]=16'hfa0f;
aud[2471]=16'hf9fa;
aud[2472]=16'hf9e5;
aud[2473]=16'hf9cf;
aud[2474]=16'hf9ba;
aud[2475]=16'hf9a5;
aud[2476]=16'hf98f;
aud[2477]=16'hf97a;
aud[2478]=16'hf965;
aud[2479]=16'hf94f;
aud[2480]=16'hf93a;
aud[2481]=16'hf925;
aud[2482]=16'hf90f;
aud[2483]=16'hf8fa;
aud[2484]=16'hf8e5;
aud[2485]=16'hf8cf;
aud[2486]=16'hf8ba;
aud[2487]=16'hf8a5;
aud[2488]=16'hf890;
aud[2489]=16'hf87a;
aud[2490]=16'hf865;
aud[2491]=16'hf850;
aud[2492]=16'hf83a;
aud[2493]=16'hf825;
aud[2494]=16'hf810;
aud[2495]=16'hf7fb;
aud[2496]=16'hf7e5;
aud[2497]=16'hf7d0;
aud[2498]=16'hf7bb;
aud[2499]=16'hf7a5;
aud[2500]=16'hf790;
aud[2501]=16'hf77b;
aud[2502]=16'hf766;
aud[2503]=16'hf750;
aud[2504]=16'hf73b;
aud[2505]=16'hf726;
aud[2506]=16'hf711;
aud[2507]=16'hf6fb;
aud[2508]=16'hf6e6;
aud[2509]=16'hf6d1;
aud[2510]=16'hf6bc;
aud[2511]=16'hf6a7;
aud[2512]=16'hf691;
aud[2513]=16'hf67c;
aud[2514]=16'hf667;
aud[2515]=16'hf652;
aud[2516]=16'hf63d;
aud[2517]=16'hf627;
aud[2518]=16'hf612;
aud[2519]=16'hf5fd;
aud[2520]=16'hf5e8;
aud[2521]=16'hf5d3;
aud[2522]=16'hf5bd;
aud[2523]=16'hf5a8;
aud[2524]=16'hf593;
aud[2525]=16'hf57e;
aud[2526]=16'hf569;
aud[2527]=16'hf554;
aud[2528]=16'hf53f;
aud[2529]=16'hf529;
aud[2530]=16'hf514;
aud[2531]=16'hf4ff;
aud[2532]=16'hf4ea;
aud[2533]=16'hf4d5;
aud[2534]=16'hf4c0;
aud[2535]=16'hf4ab;
aud[2536]=16'hf496;
aud[2537]=16'hf480;
aud[2538]=16'hf46b;
aud[2539]=16'hf456;
aud[2540]=16'hf441;
aud[2541]=16'hf42c;
aud[2542]=16'hf417;
aud[2543]=16'hf402;
aud[2544]=16'hf3ed;
aud[2545]=16'hf3d8;
aud[2546]=16'hf3c3;
aud[2547]=16'hf3ae;
aud[2548]=16'hf399;
aud[2549]=16'hf384;
aud[2550]=16'hf36f;
aud[2551]=16'hf35a;
aud[2552]=16'hf345;
aud[2553]=16'hf330;
aud[2554]=16'hf31b;
aud[2555]=16'hf306;
aud[2556]=16'hf2f1;
aud[2557]=16'hf2dc;
aud[2558]=16'hf2c7;
aud[2559]=16'hf2b2;
aud[2560]=16'hf29d;
aud[2561]=16'hf288;
aud[2562]=16'hf273;
aud[2563]=16'hf25e;
aud[2564]=16'hf249;
aud[2565]=16'hf234;
aud[2566]=16'hf21f;
aud[2567]=16'hf20a;
aud[2568]=16'hf1f5;
aud[2569]=16'hf1e0;
aud[2570]=16'hf1cb;
aud[2571]=16'hf1b6;
aud[2572]=16'hf1a1;
aud[2573]=16'hf18c;
aud[2574]=16'hf178;
aud[2575]=16'hf163;
aud[2576]=16'hf14e;
aud[2577]=16'hf139;
aud[2578]=16'hf124;
aud[2579]=16'hf10f;
aud[2580]=16'hf0fa;
aud[2581]=16'hf0e6;
aud[2582]=16'hf0d1;
aud[2583]=16'hf0bc;
aud[2584]=16'hf0a7;
aud[2585]=16'hf092;
aud[2586]=16'hf07d;
aud[2587]=16'hf069;
aud[2588]=16'hf054;
aud[2589]=16'hf03f;
aud[2590]=16'hf02a;
aud[2591]=16'hf015;
aud[2592]=16'hf001;
aud[2593]=16'hefec;
aud[2594]=16'hefd7;
aud[2595]=16'hefc2;
aud[2596]=16'hefae;
aud[2597]=16'hef99;
aud[2598]=16'hef84;
aud[2599]=16'hef70;
aud[2600]=16'hef5b;
aud[2601]=16'hef46;
aud[2602]=16'hef31;
aud[2603]=16'hef1d;
aud[2604]=16'hef08;
aud[2605]=16'heef3;
aud[2606]=16'heedf;
aud[2607]=16'heeca;
aud[2608]=16'heeb5;
aud[2609]=16'heea1;
aud[2610]=16'hee8c;
aud[2611]=16'hee77;
aud[2612]=16'hee63;
aud[2613]=16'hee4e;
aud[2614]=16'hee3a;
aud[2615]=16'hee25;
aud[2616]=16'hee10;
aud[2617]=16'hedfc;
aud[2618]=16'hede7;
aud[2619]=16'hedd3;
aud[2620]=16'hedbe;
aud[2621]=16'hedaa;
aud[2622]=16'hed95;
aud[2623]=16'hed81;
aud[2624]=16'hed6c;
aud[2625]=16'hed57;
aud[2626]=16'hed43;
aud[2627]=16'hed2e;
aud[2628]=16'hed1a;
aud[2629]=16'hed05;
aud[2630]=16'hecf1;
aud[2631]=16'hecdd;
aud[2632]=16'hecc8;
aud[2633]=16'hecb4;
aud[2634]=16'hec9f;
aud[2635]=16'hec8b;
aud[2636]=16'hec76;
aud[2637]=16'hec62;
aud[2638]=16'hec4d;
aud[2639]=16'hec39;
aud[2640]=16'hec25;
aud[2641]=16'hec10;
aud[2642]=16'hebfc;
aud[2643]=16'hebe8;
aud[2644]=16'hebd3;
aud[2645]=16'hebbf;
aud[2646]=16'hebab;
aud[2647]=16'heb96;
aud[2648]=16'heb82;
aud[2649]=16'heb6e;
aud[2650]=16'heb59;
aud[2651]=16'heb45;
aud[2652]=16'heb31;
aud[2653]=16'heb1c;
aud[2654]=16'heb08;
aud[2655]=16'heaf4;
aud[2656]=16'heae0;
aud[2657]=16'heacb;
aud[2658]=16'heab7;
aud[2659]=16'heaa3;
aud[2660]=16'hea8f;
aud[2661]=16'hea7a;
aud[2662]=16'hea66;
aud[2663]=16'hea52;
aud[2664]=16'hea3e;
aud[2665]=16'hea2a;
aud[2666]=16'hea16;
aud[2667]=16'hea01;
aud[2668]=16'he9ed;
aud[2669]=16'he9d9;
aud[2670]=16'he9c5;
aud[2671]=16'he9b1;
aud[2672]=16'he99d;
aud[2673]=16'he989;
aud[2674]=16'he975;
aud[2675]=16'he961;
aud[2676]=16'he94d;
aud[2677]=16'he939;
aud[2678]=16'he925;
aud[2679]=16'he910;
aud[2680]=16'he8fc;
aud[2681]=16'he8e8;
aud[2682]=16'he8d4;
aud[2683]=16'he8c0;
aud[2684]=16'he8ad;
aud[2685]=16'he899;
aud[2686]=16'he885;
aud[2687]=16'he871;
aud[2688]=16'he85d;
aud[2689]=16'he849;
aud[2690]=16'he835;
aud[2691]=16'he821;
aud[2692]=16'he80d;
aud[2693]=16'he7f9;
aud[2694]=16'he7e5;
aud[2695]=16'he7d1;
aud[2696]=16'he7be;
aud[2697]=16'he7aa;
aud[2698]=16'he796;
aud[2699]=16'he782;
aud[2700]=16'he76e;
aud[2701]=16'he75b;
aud[2702]=16'he747;
aud[2703]=16'he733;
aud[2704]=16'he71f;
aud[2705]=16'he70b;
aud[2706]=16'he6f8;
aud[2707]=16'he6e4;
aud[2708]=16'he6d0;
aud[2709]=16'he6bd;
aud[2710]=16'he6a9;
aud[2711]=16'he695;
aud[2712]=16'he681;
aud[2713]=16'he66e;
aud[2714]=16'he65a;
aud[2715]=16'he646;
aud[2716]=16'he633;
aud[2717]=16'he61f;
aud[2718]=16'he60c;
aud[2719]=16'he5f8;
aud[2720]=16'he5e4;
aud[2721]=16'he5d1;
aud[2722]=16'he5bd;
aud[2723]=16'he5aa;
aud[2724]=16'he596;
aud[2725]=16'he583;
aud[2726]=16'he56f;
aud[2727]=16'he55c;
aud[2728]=16'he548;
aud[2729]=16'he535;
aud[2730]=16'he521;
aud[2731]=16'he50e;
aud[2732]=16'he4fa;
aud[2733]=16'he4e7;
aud[2734]=16'he4d3;
aud[2735]=16'he4c0;
aud[2736]=16'he4ad;
aud[2737]=16'he499;
aud[2738]=16'he486;
aud[2739]=16'he473;
aud[2740]=16'he45f;
aud[2741]=16'he44c;
aud[2742]=16'he438;
aud[2743]=16'he425;
aud[2744]=16'he412;
aud[2745]=16'he3ff;
aud[2746]=16'he3eb;
aud[2747]=16'he3d8;
aud[2748]=16'he3c5;
aud[2749]=16'he3b2;
aud[2750]=16'he39e;
aud[2751]=16'he38b;
aud[2752]=16'he378;
aud[2753]=16'he365;
aud[2754]=16'he352;
aud[2755]=16'he33e;
aud[2756]=16'he32b;
aud[2757]=16'he318;
aud[2758]=16'he305;
aud[2759]=16'he2f2;
aud[2760]=16'he2df;
aud[2761]=16'he2cc;
aud[2762]=16'he2b9;
aud[2763]=16'he2a5;
aud[2764]=16'he292;
aud[2765]=16'he27f;
aud[2766]=16'he26c;
aud[2767]=16'he259;
aud[2768]=16'he246;
aud[2769]=16'he233;
aud[2770]=16'he220;
aud[2771]=16'he20d;
aud[2772]=16'he1fa;
aud[2773]=16'he1e8;
aud[2774]=16'he1d5;
aud[2775]=16'he1c2;
aud[2776]=16'he1af;
aud[2777]=16'he19c;
aud[2778]=16'he189;
aud[2779]=16'he176;
aud[2780]=16'he163;
aud[2781]=16'he151;
aud[2782]=16'he13e;
aud[2783]=16'he12b;
aud[2784]=16'he118;
aud[2785]=16'he105;
aud[2786]=16'he0f3;
aud[2787]=16'he0e0;
aud[2788]=16'he0cd;
aud[2789]=16'he0ba;
aud[2790]=16'he0a8;
aud[2791]=16'he095;
aud[2792]=16'he082;
aud[2793]=16'he070;
aud[2794]=16'he05d;
aud[2795]=16'he04a;
aud[2796]=16'he038;
aud[2797]=16'he025;
aud[2798]=16'he013;
aud[2799]=16'he000;
aud[2800]=16'hdfed;
aud[2801]=16'hdfdb;
aud[2802]=16'hdfc8;
aud[2803]=16'hdfb6;
aud[2804]=16'hdfa3;
aud[2805]=16'hdf91;
aud[2806]=16'hdf7e;
aud[2807]=16'hdf6c;
aud[2808]=16'hdf59;
aud[2809]=16'hdf47;
aud[2810]=16'hdf35;
aud[2811]=16'hdf22;
aud[2812]=16'hdf10;
aud[2813]=16'hdefd;
aud[2814]=16'hdeeb;
aud[2815]=16'hded9;
aud[2816]=16'hdec6;
aud[2817]=16'hdeb4;
aud[2818]=16'hdea2;
aud[2819]=16'hde8f;
aud[2820]=16'hde7d;
aud[2821]=16'hde6b;
aud[2822]=16'hde59;
aud[2823]=16'hde46;
aud[2824]=16'hde34;
aud[2825]=16'hde22;
aud[2826]=16'hde10;
aud[2827]=16'hddfe;
aud[2828]=16'hddeb;
aud[2829]=16'hddd9;
aud[2830]=16'hddc7;
aud[2831]=16'hddb5;
aud[2832]=16'hdda3;
aud[2833]=16'hdd91;
aud[2834]=16'hdd7f;
aud[2835]=16'hdd6d;
aud[2836]=16'hdd5b;
aud[2837]=16'hdd49;
aud[2838]=16'hdd37;
aud[2839]=16'hdd25;
aud[2840]=16'hdd13;
aud[2841]=16'hdd01;
aud[2842]=16'hdcef;
aud[2843]=16'hdcdd;
aud[2844]=16'hdccb;
aud[2845]=16'hdcb9;
aud[2846]=16'hdca7;
aud[2847]=16'hdc95;
aud[2848]=16'hdc83;
aud[2849]=16'hdc72;
aud[2850]=16'hdc60;
aud[2851]=16'hdc4e;
aud[2852]=16'hdc3c;
aud[2853]=16'hdc2a;
aud[2854]=16'hdc19;
aud[2855]=16'hdc07;
aud[2856]=16'hdbf5;
aud[2857]=16'hdbe3;
aud[2858]=16'hdbd2;
aud[2859]=16'hdbc0;
aud[2860]=16'hdbae;
aud[2861]=16'hdb9d;
aud[2862]=16'hdb8b;
aud[2863]=16'hdb79;
aud[2864]=16'hdb68;
aud[2865]=16'hdb56;
aud[2866]=16'hdb45;
aud[2867]=16'hdb33;
aud[2868]=16'hdb22;
aud[2869]=16'hdb10;
aud[2870]=16'hdaff;
aud[2871]=16'hdaed;
aud[2872]=16'hdadc;
aud[2873]=16'hdaca;
aud[2874]=16'hdab9;
aud[2875]=16'hdaa7;
aud[2876]=16'hda96;
aud[2877]=16'hda84;
aud[2878]=16'hda73;
aud[2879]=16'hda62;
aud[2880]=16'hda50;
aud[2881]=16'hda3f;
aud[2882]=16'hda2e;
aud[2883]=16'hda1c;
aud[2884]=16'hda0b;
aud[2885]=16'hd9fa;
aud[2886]=16'hd9e9;
aud[2887]=16'hd9d7;
aud[2888]=16'hd9c6;
aud[2889]=16'hd9b5;
aud[2890]=16'hd9a4;
aud[2891]=16'hd993;
aud[2892]=16'hd982;
aud[2893]=16'hd970;
aud[2894]=16'hd95f;
aud[2895]=16'hd94e;
aud[2896]=16'hd93d;
aud[2897]=16'hd92c;
aud[2898]=16'hd91b;
aud[2899]=16'hd90a;
aud[2900]=16'hd8f9;
aud[2901]=16'hd8e8;
aud[2902]=16'hd8d7;
aud[2903]=16'hd8c6;
aud[2904]=16'hd8b5;
aud[2905]=16'hd8a4;
aud[2906]=16'hd893;
aud[2907]=16'hd882;
aud[2908]=16'hd872;
aud[2909]=16'hd861;
aud[2910]=16'hd850;
aud[2911]=16'hd83f;
aud[2912]=16'hd82e;
aud[2913]=16'hd81e;
aud[2914]=16'hd80d;
aud[2915]=16'hd7fc;
aud[2916]=16'hd7eb;
aud[2917]=16'hd7db;
aud[2918]=16'hd7ca;
aud[2919]=16'hd7b9;
aud[2920]=16'hd7a9;
aud[2921]=16'hd798;
aud[2922]=16'hd787;
aud[2923]=16'hd777;
aud[2924]=16'hd766;
aud[2925]=16'hd756;
aud[2926]=16'hd745;
aud[2927]=16'hd734;
aud[2928]=16'hd724;
aud[2929]=16'hd713;
aud[2930]=16'hd703;
aud[2931]=16'hd6f2;
aud[2932]=16'hd6e2;
aud[2933]=16'hd6d2;
aud[2934]=16'hd6c1;
aud[2935]=16'hd6b1;
aud[2936]=16'hd6a0;
aud[2937]=16'hd690;
aud[2938]=16'hd680;
aud[2939]=16'hd66f;
aud[2940]=16'hd65f;
aud[2941]=16'hd64f;
aud[2942]=16'hd63f;
aud[2943]=16'hd62e;
aud[2944]=16'hd61e;
aud[2945]=16'hd60e;
aud[2946]=16'hd5fe;
aud[2947]=16'hd5ee;
aud[2948]=16'hd5dd;
aud[2949]=16'hd5cd;
aud[2950]=16'hd5bd;
aud[2951]=16'hd5ad;
aud[2952]=16'hd59d;
aud[2953]=16'hd58d;
aud[2954]=16'hd57d;
aud[2955]=16'hd56d;
aud[2956]=16'hd55d;
aud[2957]=16'hd54d;
aud[2958]=16'hd53d;
aud[2959]=16'hd52d;
aud[2960]=16'hd51d;
aud[2961]=16'hd50d;
aud[2962]=16'hd4fd;
aud[2963]=16'hd4ed;
aud[2964]=16'hd4de;
aud[2965]=16'hd4ce;
aud[2966]=16'hd4be;
aud[2967]=16'hd4ae;
aud[2968]=16'hd49e;
aud[2969]=16'hd48f;
aud[2970]=16'hd47f;
aud[2971]=16'hd46f;
aud[2972]=16'hd45f;
aud[2973]=16'hd450;
aud[2974]=16'hd440;
aud[2975]=16'hd430;
aud[2976]=16'hd421;
aud[2977]=16'hd411;
aud[2978]=16'hd402;
aud[2979]=16'hd3f2;
aud[2980]=16'hd3e2;
aud[2981]=16'hd3d3;
aud[2982]=16'hd3c3;
aud[2983]=16'hd3b4;
aud[2984]=16'hd3a4;
aud[2985]=16'hd395;
aud[2986]=16'hd386;
aud[2987]=16'hd376;
aud[2988]=16'hd367;
aud[2989]=16'hd357;
aud[2990]=16'hd348;
aud[2991]=16'hd339;
aud[2992]=16'hd329;
aud[2993]=16'hd31a;
aud[2994]=16'hd30b;
aud[2995]=16'hd2fc;
aud[2996]=16'hd2ec;
aud[2997]=16'hd2dd;
aud[2998]=16'hd2ce;
aud[2999]=16'hd2bf;
aud[3000]=16'hd2b0;
aud[3001]=16'hd2a0;
aud[3002]=16'hd291;
aud[3003]=16'hd282;
aud[3004]=16'hd273;
aud[3005]=16'hd264;
aud[3006]=16'hd255;
aud[3007]=16'hd246;
aud[3008]=16'hd237;
aud[3009]=16'hd228;
aud[3010]=16'hd219;
aud[3011]=16'hd20a;
aud[3012]=16'hd1fb;
aud[3013]=16'hd1ec;
aud[3014]=16'hd1de;
aud[3015]=16'hd1cf;
aud[3016]=16'hd1c0;
aud[3017]=16'hd1b1;
aud[3018]=16'hd1a2;
aud[3019]=16'hd193;
aud[3020]=16'hd185;
aud[3021]=16'hd176;
aud[3022]=16'hd167;
aud[3023]=16'hd159;
aud[3024]=16'hd14a;
aud[3025]=16'hd13b;
aud[3026]=16'hd12d;
aud[3027]=16'hd11e;
aud[3028]=16'hd10f;
aud[3029]=16'hd101;
aud[3030]=16'hd0f2;
aud[3031]=16'hd0e4;
aud[3032]=16'hd0d5;
aud[3033]=16'hd0c7;
aud[3034]=16'hd0b8;
aud[3035]=16'hd0aa;
aud[3036]=16'hd09b;
aud[3037]=16'hd08d;
aud[3038]=16'hd07f;
aud[3039]=16'hd070;
aud[3040]=16'hd062;
aud[3041]=16'hd054;
aud[3042]=16'hd045;
aud[3043]=16'hd037;
aud[3044]=16'hd029;
aud[3045]=16'hd01b;
aud[3046]=16'hd00c;
aud[3047]=16'hcffe;
aud[3048]=16'hcff0;
aud[3049]=16'hcfe2;
aud[3050]=16'hcfd4;
aud[3051]=16'hcfc6;
aud[3052]=16'hcfb8;
aud[3053]=16'hcfa9;
aud[3054]=16'hcf9b;
aud[3055]=16'hcf8d;
aud[3056]=16'hcf7f;
aud[3057]=16'hcf71;
aud[3058]=16'hcf63;
aud[3059]=16'hcf56;
aud[3060]=16'hcf48;
aud[3061]=16'hcf3a;
aud[3062]=16'hcf2c;
aud[3063]=16'hcf1e;
aud[3064]=16'hcf10;
aud[3065]=16'hcf02;
aud[3066]=16'hcef5;
aud[3067]=16'hcee7;
aud[3068]=16'hced9;
aud[3069]=16'hcecb;
aud[3070]=16'hcebe;
aud[3071]=16'hceb0;
aud[3072]=16'hcea2;
aud[3073]=16'hce95;
aud[3074]=16'hce87;
aud[3075]=16'hce79;
aud[3076]=16'hce6c;
aud[3077]=16'hce5e;
aud[3078]=16'hce51;
aud[3079]=16'hce43;
aud[3080]=16'hce36;
aud[3081]=16'hce28;
aud[3082]=16'hce1b;
aud[3083]=16'hce0d;
aud[3084]=16'hce00;
aud[3085]=16'hcdf3;
aud[3086]=16'hcde5;
aud[3087]=16'hcdd8;
aud[3088]=16'hcdcb;
aud[3089]=16'hcdbd;
aud[3090]=16'hcdb0;
aud[3091]=16'hcda3;
aud[3092]=16'hcd96;
aud[3093]=16'hcd88;
aud[3094]=16'hcd7b;
aud[3095]=16'hcd6e;
aud[3096]=16'hcd61;
aud[3097]=16'hcd54;
aud[3098]=16'hcd47;
aud[3099]=16'hcd3a;
aud[3100]=16'hcd2d;
aud[3101]=16'hcd20;
aud[3102]=16'hcd13;
aud[3103]=16'hcd06;
aud[3104]=16'hccf9;
aud[3105]=16'hccec;
aud[3106]=16'hccdf;
aud[3107]=16'hccd2;
aud[3108]=16'hccc5;
aud[3109]=16'hccb8;
aud[3110]=16'hccab;
aud[3111]=16'hcc9f;
aud[3112]=16'hcc92;
aud[3113]=16'hcc85;
aud[3114]=16'hcc78;
aud[3115]=16'hcc6c;
aud[3116]=16'hcc5f;
aud[3117]=16'hcc52;
aud[3118]=16'hcc46;
aud[3119]=16'hcc39;
aud[3120]=16'hcc2c;
aud[3121]=16'hcc20;
aud[3122]=16'hcc13;
aud[3123]=16'hcc07;
aud[3124]=16'hcbfa;
aud[3125]=16'hcbee;
aud[3126]=16'hcbe1;
aud[3127]=16'hcbd5;
aud[3128]=16'hcbc9;
aud[3129]=16'hcbbc;
aud[3130]=16'hcbb0;
aud[3131]=16'hcba3;
aud[3132]=16'hcb97;
aud[3133]=16'hcb8b;
aud[3134]=16'hcb7f;
aud[3135]=16'hcb72;
aud[3136]=16'hcb66;
aud[3137]=16'hcb5a;
aud[3138]=16'hcb4e;
aud[3139]=16'hcb42;
aud[3140]=16'hcb35;
aud[3141]=16'hcb29;
aud[3142]=16'hcb1d;
aud[3143]=16'hcb11;
aud[3144]=16'hcb05;
aud[3145]=16'hcaf9;
aud[3146]=16'hcaed;
aud[3147]=16'hcae1;
aud[3148]=16'hcad5;
aud[3149]=16'hcac9;
aud[3150]=16'hcabd;
aud[3151]=16'hcab1;
aud[3152]=16'hcaa6;
aud[3153]=16'hca9a;
aud[3154]=16'hca8e;
aud[3155]=16'hca82;
aud[3156]=16'hca76;
aud[3157]=16'hca6b;
aud[3158]=16'hca5f;
aud[3159]=16'hca53;
aud[3160]=16'hca48;
aud[3161]=16'hca3c;
aud[3162]=16'hca30;
aud[3163]=16'hca25;
aud[3164]=16'hca19;
aud[3165]=16'hca0e;
aud[3166]=16'hca02;
aud[3167]=16'hc9f7;
aud[3168]=16'hc9eb;
aud[3169]=16'hc9e0;
aud[3170]=16'hc9d4;
aud[3171]=16'hc9c9;
aud[3172]=16'hc9bd;
aud[3173]=16'hc9b2;
aud[3174]=16'hc9a7;
aud[3175]=16'hc99b;
aud[3176]=16'hc990;
aud[3177]=16'hc985;
aud[3178]=16'hc97a;
aud[3179]=16'hc96e;
aud[3180]=16'hc963;
aud[3181]=16'hc958;
aud[3182]=16'hc94d;
aud[3183]=16'hc942;
aud[3184]=16'hc937;
aud[3185]=16'hc92c;
aud[3186]=16'hc920;
aud[3187]=16'hc915;
aud[3188]=16'hc90a;
aud[3189]=16'hc8ff;
aud[3190]=16'hc8f5;
aud[3191]=16'hc8ea;
aud[3192]=16'hc8df;
aud[3193]=16'hc8d4;
aud[3194]=16'hc8c9;
aud[3195]=16'hc8be;
aud[3196]=16'hc8b3;
aud[3197]=16'hc8a9;
aud[3198]=16'hc89e;
aud[3199]=16'hc893;
aud[3200]=16'hc888;
aud[3201]=16'hc87e;
aud[3202]=16'hc873;
aud[3203]=16'hc868;
aud[3204]=16'hc85e;
aud[3205]=16'hc853;
aud[3206]=16'hc849;
aud[3207]=16'hc83e;
aud[3208]=16'hc834;
aud[3209]=16'hc829;
aud[3210]=16'hc81f;
aud[3211]=16'hc814;
aud[3212]=16'hc80a;
aud[3213]=16'hc7ff;
aud[3214]=16'hc7f5;
aud[3215]=16'hc7eb;
aud[3216]=16'hc7e0;
aud[3217]=16'hc7d6;
aud[3218]=16'hc7cc;
aud[3219]=16'hc7c1;
aud[3220]=16'hc7b7;
aud[3221]=16'hc7ad;
aud[3222]=16'hc7a3;
aud[3223]=16'hc799;
aud[3224]=16'hc78f;
aud[3225]=16'hc785;
aud[3226]=16'hc77a;
aud[3227]=16'hc770;
aud[3228]=16'hc766;
aud[3229]=16'hc75c;
aud[3230]=16'hc752;
aud[3231]=16'hc748;
aud[3232]=16'hc73f;
aud[3233]=16'hc735;
aud[3234]=16'hc72b;
aud[3235]=16'hc721;
aud[3236]=16'hc717;
aud[3237]=16'hc70d;
aud[3238]=16'hc703;
aud[3239]=16'hc6fa;
aud[3240]=16'hc6f0;
aud[3241]=16'hc6e6;
aud[3242]=16'hc6dd;
aud[3243]=16'hc6d3;
aud[3244]=16'hc6c9;
aud[3245]=16'hc6c0;
aud[3246]=16'hc6b6;
aud[3247]=16'hc6ad;
aud[3248]=16'hc6a3;
aud[3249]=16'hc69a;
aud[3250]=16'hc690;
aud[3251]=16'hc687;
aud[3252]=16'hc67d;
aud[3253]=16'hc674;
aud[3254]=16'hc66b;
aud[3255]=16'hc661;
aud[3256]=16'hc658;
aud[3257]=16'hc64f;
aud[3258]=16'hc645;
aud[3259]=16'hc63c;
aud[3260]=16'hc633;
aud[3261]=16'hc62a;
aud[3262]=16'hc620;
aud[3263]=16'hc617;
aud[3264]=16'hc60e;
aud[3265]=16'hc605;
aud[3266]=16'hc5fc;
aud[3267]=16'hc5f3;
aud[3268]=16'hc5ea;
aud[3269]=16'hc5e1;
aud[3270]=16'hc5d8;
aud[3271]=16'hc5cf;
aud[3272]=16'hc5c6;
aud[3273]=16'hc5bd;
aud[3274]=16'hc5b4;
aud[3275]=16'hc5ac;
aud[3276]=16'hc5a3;
aud[3277]=16'hc59a;
aud[3278]=16'hc591;
aud[3279]=16'hc588;
aud[3280]=16'hc580;
aud[3281]=16'hc577;
aud[3282]=16'hc56e;
aud[3283]=16'hc566;
aud[3284]=16'hc55d;
aud[3285]=16'hc555;
aud[3286]=16'hc54c;
aud[3287]=16'hc544;
aud[3288]=16'hc53b;
aud[3289]=16'hc533;
aud[3290]=16'hc52a;
aud[3291]=16'hc522;
aud[3292]=16'hc519;
aud[3293]=16'hc511;
aud[3294]=16'hc509;
aud[3295]=16'hc500;
aud[3296]=16'hc4f8;
aud[3297]=16'hc4f0;
aud[3298]=16'hc4e7;
aud[3299]=16'hc4df;
aud[3300]=16'hc4d7;
aud[3301]=16'hc4cf;
aud[3302]=16'hc4c7;
aud[3303]=16'hc4bf;
aud[3304]=16'hc4b6;
aud[3305]=16'hc4ae;
aud[3306]=16'hc4a6;
aud[3307]=16'hc49e;
aud[3308]=16'hc496;
aud[3309]=16'hc48e;
aud[3310]=16'hc486;
aud[3311]=16'hc47f;
aud[3312]=16'hc477;
aud[3313]=16'hc46f;
aud[3314]=16'hc467;
aud[3315]=16'hc45f;
aud[3316]=16'hc457;
aud[3317]=16'hc450;
aud[3318]=16'hc448;
aud[3319]=16'hc440;
aud[3320]=16'hc439;
aud[3321]=16'hc431;
aud[3322]=16'hc429;
aud[3323]=16'hc422;
aud[3324]=16'hc41a;
aud[3325]=16'hc413;
aud[3326]=16'hc40b;
aud[3327]=16'hc404;
aud[3328]=16'hc3fc;
aud[3329]=16'hc3f5;
aud[3330]=16'hc3ed;
aud[3331]=16'hc3e6;
aud[3332]=16'hc3df;
aud[3333]=16'hc3d7;
aud[3334]=16'hc3d0;
aud[3335]=16'hc3c9;
aud[3336]=16'hc3c1;
aud[3337]=16'hc3ba;
aud[3338]=16'hc3b3;
aud[3339]=16'hc3ac;
aud[3340]=16'hc3a5;
aud[3341]=16'hc39d;
aud[3342]=16'hc396;
aud[3343]=16'hc38f;
aud[3344]=16'hc388;
aud[3345]=16'hc381;
aud[3346]=16'hc37a;
aud[3347]=16'hc373;
aud[3348]=16'hc36c;
aud[3349]=16'hc365;
aud[3350]=16'hc35f;
aud[3351]=16'hc358;
aud[3352]=16'hc351;
aud[3353]=16'hc34a;
aud[3354]=16'hc343;
aud[3355]=16'hc33d;
aud[3356]=16'hc336;
aud[3357]=16'hc32f;
aud[3358]=16'hc329;
aud[3359]=16'hc322;
aud[3360]=16'hc31b;
aud[3361]=16'hc315;
aud[3362]=16'hc30e;
aud[3363]=16'hc308;
aud[3364]=16'hc301;
aud[3365]=16'hc2fb;
aud[3366]=16'hc2f4;
aud[3367]=16'hc2ee;
aud[3368]=16'hc2e7;
aud[3369]=16'hc2e1;
aud[3370]=16'hc2db;
aud[3371]=16'hc2d4;
aud[3372]=16'hc2ce;
aud[3373]=16'hc2c8;
aud[3374]=16'hc2c1;
aud[3375]=16'hc2bb;
aud[3376]=16'hc2b5;
aud[3377]=16'hc2af;
aud[3378]=16'hc2a9;
aud[3379]=16'hc2a3;
aud[3380]=16'hc29d;
aud[3381]=16'hc297;
aud[3382]=16'hc291;
aud[3383]=16'hc28b;
aud[3384]=16'hc285;
aud[3385]=16'hc27f;
aud[3386]=16'hc279;
aud[3387]=16'hc273;
aud[3388]=16'hc26d;
aud[3389]=16'hc267;
aud[3390]=16'hc261;
aud[3391]=16'hc25c;
aud[3392]=16'hc256;
aud[3393]=16'hc250;
aud[3394]=16'hc24a;
aud[3395]=16'hc245;
aud[3396]=16'hc23f;
aud[3397]=16'hc239;
aud[3398]=16'hc234;
aud[3399]=16'hc22e;
aud[3400]=16'hc229;
aud[3401]=16'hc223;
aud[3402]=16'hc21e;
aud[3403]=16'hc218;
aud[3404]=16'hc213;
aud[3405]=16'hc20d;
aud[3406]=16'hc208;
aud[3407]=16'hc203;
aud[3408]=16'hc1fd;
aud[3409]=16'hc1f8;
aud[3410]=16'hc1f3;
aud[3411]=16'hc1ee;
aud[3412]=16'hc1e8;
aud[3413]=16'hc1e3;
aud[3414]=16'hc1de;
aud[3415]=16'hc1d9;
aud[3416]=16'hc1d4;
aud[3417]=16'hc1cf;
aud[3418]=16'hc1ca;
aud[3419]=16'hc1c5;
aud[3420]=16'hc1c0;
aud[3421]=16'hc1bb;
aud[3422]=16'hc1b6;
aud[3423]=16'hc1b1;
aud[3424]=16'hc1ac;
aud[3425]=16'hc1a7;
aud[3426]=16'hc1a2;
aud[3427]=16'hc19e;
aud[3428]=16'hc199;
aud[3429]=16'hc194;
aud[3430]=16'hc18f;
aud[3431]=16'hc18b;
aud[3432]=16'hc186;
aud[3433]=16'hc181;
aud[3434]=16'hc17d;
aud[3435]=16'hc178;
aud[3436]=16'hc174;
aud[3437]=16'hc16f;
aud[3438]=16'hc16b;
aud[3439]=16'hc166;
aud[3440]=16'hc162;
aud[3441]=16'hc15d;
aud[3442]=16'hc159;
aud[3443]=16'hc154;
aud[3444]=16'hc150;
aud[3445]=16'hc14c;
aud[3446]=16'hc147;
aud[3447]=16'hc143;
aud[3448]=16'hc13f;
aud[3449]=16'hc13b;
aud[3450]=16'hc137;
aud[3451]=16'hc133;
aud[3452]=16'hc12e;
aud[3453]=16'hc12a;
aud[3454]=16'hc126;
aud[3455]=16'hc122;
aud[3456]=16'hc11e;
aud[3457]=16'hc11a;
aud[3458]=16'hc116;
aud[3459]=16'hc112;
aud[3460]=16'hc10e;
aud[3461]=16'hc10b;
aud[3462]=16'hc107;
aud[3463]=16'hc103;
aud[3464]=16'hc0ff;
aud[3465]=16'hc0fb;
aud[3466]=16'hc0f8;
aud[3467]=16'hc0f4;
aud[3468]=16'hc0f0;
aud[3469]=16'hc0ed;
aud[3470]=16'hc0e9;
aud[3471]=16'hc0e5;
aud[3472]=16'hc0e2;
aud[3473]=16'hc0de;
aud[3474]=16'hc0db;
aud[3475]=16'hc0d7;
aud[3476]=16'hc0d4;
aud[3477]=16'hc0d0;
aud[3478]=16'hc0cd;
aud[3479]=16'hc0ca;
aud[3480]=16'hc0c6;
aud[3481]=16'hc0c3;
aud[3482]=16'hc0c0;
aud[3483]=16'hc0bd;
aud[3484]=16'hc0b9;
aud[3485]=16'hc0b6;
aud[3486]=16'hc0b3;
aud[3487]=16'hc0b0;
aud[3488]=16'hc0ad;
aud[3489]=16'hc0aa;
aud[3490]=16'hc0a6;
aud[3491]=16'hc0a3;
aud[3492]=16'hc0a0;
aud[3493]=16'hc09d;
aud[3494]=16'hc09b;
aud[3495]=16'hc098;
aud[3496]=16'hc095;
aud[3497]=16'hc092;
aud[3498]=16'hc08f;
aud[3499]=16'hc08c;
aud[3500]=16'hc089;
aud[3501]=16'hc087;
aud[3502]=16'hc084;
aud[3503]=16'hc081;
aud[3504]=16'hc07f;
aud[3505]=16'hc07c;
aud[3506]=16'hc079;
aud[3507]=16'hc077;
aud[3508]=16'hc074;
aud[3509]=16'hc072;
aud[3510]=16'hc06f;
aud[3511]=16'hc06d;
aud[3512]=16'hc06a;
aud[3513]=16'hc068;
aud[3514]=16'hc065;
aud[3515]=16'hc063;
aud[3516]=16'hc061;
aud[3517]=16'hc05e;
aud[3518]=16'hc05c;
aud[3519]=16'hc05a;
aud[3520]=16'hc058;
aud[3521]=16'hc055;
aud[3522]=16'hc053;
aud[3523]=16'hc051;
aud[3524]=16'hc04f;
aud[3525]=16'hc04d;
aud[3526]=16'hc04b;
aud[3527]=16'hc049;
aud[3528]=16'hc047;
aud[3529]=16'hc045;
aud[3530]=16'hc043;
aud[3531]=16'hc041;
aud[3532]=16'hc03f;
aud[3533]=16'hc03d;
aud[3534]=16'hc03b;
aud[3535]=16'hc039;
aud[3536]=16'hc038;
aud[3537]=16'hc036;
aud[3538]=16'hc034;
aud[3539]=16'hc033;
aud[3540]=16'hc031;
aud[3541]=16'hc02f;
aud[3542]=16'hc02e;
aud[3543]=16'hc02c;
aud[3544]=16'hc02a;
aud[3545]=16'hc029;
aud[3546]=16'hc027;
aud[3547]=16'hc026;
aud[3548]=16'hc024;
aud[3549]=16'hc023;
aud[3550]=16'hc022;
aud[3551]=16'hc020;
aud[3552]=16'hc01f;
aud[3553]=16'hc01e;
aud[3554]=16'hc01c;
aud[3555]=16'hc01b;
aud[3556]=16'hc01a;
aud[3557]=16'hc019;
aud[3558]=16'hc018;
aud[3559]=16'hc016;
aud[3560]=16'hc015;
aud[3561]=16'hc014;
aud[3562]=16'hc013;
aud[3563]=16'hc012;
aud[3564]=16'hc011;
aud[3565]=16'hc010;
aud[3566]=16'hc00f;
aud[3567]=16'hc00e;
aud[3568]=16'hc00d;
aud[3569]=16'hc00d;
aud[3570]=16'hc00c;
aud[3571]=16'hc00b;
aud[3572]=16'hc00a;
aud[3573]=16'hc009;
aud[3574]=16'hc009;
aud[3575]=16'hc008;
aud[3576]=16'hc007;
aud[3577]=16'hc007;
aud[3578]=16'hc006;
aud[3579]=16'hc006;
aud[3580]=16'hc005;
aud[3581]=16'hc005;
aud[3582]=16'hc004;
aud[3583]=16'hc004;
aud[3584]=16'hc003;
aud[3585]=16'hc003;
aud[3586]=16'hc002;
aud[3587]=16'hc002;
aud[3588]=16'hc002;
aud[3589]=16'hc001;
aud[3590]=16'hc001;
aud[3591]=16'hc001;
aud[3592]=16'hc001;
aud[3593]=16'hc001;
aud[3594]=16'hc000;
aud[3595]=16'hc000;
aud[3596]=16'hc000;
aud[3597]=16'hc000;
aud[3598]=16'hc000;
aud[3599]=16'hc000;
aud[3600]=16'hc000;
aud[3601]=16'hc000;
aud[3602]=16'hc000;
aud[3603]=16'hc000;
aud[3604]=16'hc000;
aud[3605]=16'hc001;
aud[3606]=16'hc001;
aud[3607]=16'hc001;
aud[3608]=16'hc001;
aud[3609]=16'hc001;
aud[3610]=16'hc002;
aud[3611]=16'hc002;
aud[3612]=16'hc002;
aud[3613]=16'hc003;
aud[3614]=16'hc003;
aud[3615]=16'hc004;
aud[3616]=16'hc004;
aud[3617]=16'hc005;
aud[3618]=16'hc005;
aud[3619]=16'hc006;
aud[3620]=16'hc006;
aud[3621]=16'hc007;
aud[3622]=16'hc007;
aud[3623]=16'hc008;
aud[3624]=16'hc009;
aud[3625]=16'hc009;
aud[3626]=16'hc00a;
aud[3627]=16'hc00b;
aud[3628]=16'hc00c;
aud[3629]=16'hc00d;
aud[3630]=16'hc00d;
aud[3631]=16'hc00e;
aud[3632]=16'hc00f;
aud[3633]=16'hc010;
aud[3634]=16'hc011;
aud[3635]=16'hc012;
aud[3636]=16'hc013;
aud[3637]=16'hc014;
aud[3638]=16'hc015;
aud[3639]=16'hc016;
aud[3640]=16'hc018;
aud[3641]=16'hc019;
aud[3642]=16'hc01a;
aud[3643]=16'hc01b;
aud[3644]=16'hc01c;
aud[3645]=16'hc01e;
aud[3646]=16'hc01f;
aud[3647]=16'hc020;
aud[3648]=16'hc022;
aud[3649]=16'hc023;
aud[3650]=16'hc024;
aud[3651]=16'hc026;
aud[3652]=16'hc027;
aud[3653]=16'hc029;
aud[3654]=16'hc02a;
aud[3655]=16'hc02c;
aud[3656]=16'hc02e;
aud[3657]=16'hc02f;
aud[3658]=16'hc031;
aud[3659]=16'hc033;
aud[3660]=16'hc034;
aud[3661]=16'hc036;
aud[3662]=16'hc038;
aud[3663]=16'hc039;
aud[3664]=16'hc03b;
aud[3665]=16'hc03d;
aud[3666]=16'hc03f;
aud[3667]=16'hc041;
aud[3668]=16'hc043;
aud[3669]=16'hc045;
aud[3670]=16'hc047;
aud[3671]=16'hc049;
aud[3672]=16'hc04b;
aud[3673]=16'hc04d;
aud[3674]=16'hc04f;
aud[3675]=16'hc051;
aud[3676]=16'hc053;
aud[3677]=16'hc055;
aud[3678]=16'hc058;
aud[3679]=16'hc05a;
aud[3680]=16'hc05c;
aud[3681]=16'hc05e;
aud[3682]=16'hc061;
aud[3683]=16'hc063;
aud[3684]=16'hc065;
aud[3685]=16'hc068;
aud[3686]=16'hc06a;
aud[3687]=16'hc06d;
aud[3688]=16'hc06f;
aud[3689]=16'hc072;
aud[3690]=16'hc074;
aud[3691]=16'hc077;
aud[3692]=16'hc079;
aud[3693]=16'hc07c;
aud[3694]=16'hc07f;
aud[3695]=16'hc081;
aud[3696]=16'hc084;
aud[3697]=16'hc087;
aud[3698]=16'hc089;
aud[3699]=16'hc08c;
aud[3700]=16'hc08f;
aud[3701]=16'hc092;
aud[3702]=16'hc095;
aud[3703]=16'hc098;
aud[3704]=16'hc09b;
aud[3705]=16'hc09d;
aud[3706]=16'hc0a0;
aud[3707]=16'hc0a3;
aud[3708]=16'hc0a6;
aud[3709]=16'hc0aa;
aud[3710]=16'hc0ad;
aud[3711]=16'hc0b0;
aud[3712]=16'hc0b3;
aud[3713]=16'hc0b6;
aud[3714]=16'hc0b9;
aud[3715]=16'hc0bd;
aud[3716]=16'hc0c0;
aud[3717]=16'hc0c3;
aud[3718]=16'hc0c6;
aud[3719]=16'hc0ca;
aud[3720]=16'hc0cd;
aud[3721]=16'hc0d0;
aud[3722]=16'hc0d4;
aud[3723]=16'hc0d7;
aud[3724]=16'hc0db;
aud[3725]=16'hc0de;
aud[3726]=16'hc0e2;
aud[3727]=16'hc0e5;
aud[3728]=16'hc0e9;
aud[3729]=16'hc0ed;
aud[3730]=16'hc0f0;
aud[3731]=16'hc0f4;
aud[3732]=16'hc0f8;
aud[3733]=16'hc0fb;
aud[3734]=16'hc0ff;
aud[3735]=16'hc103;
aud[3736]=16'hc107;
aud[3737]=16'hc10b;
aud[3738]=16'hc10e;
aud[3739]=16'hc112;
aud[3740]=16'hc116;
aud[3741]=16'hc11a;
aud[3742]=16'hc11e;
aud[3743]=16'hc122;
aud[3744]=16'hc126;
aud[3745]=16'hc12a;
aud[3746]=16'hc12e;
aud[3747]=16'hc133;
aud[3748]=16'hc137;
aud[3749]=16'hc13b;
aud[3750]=16'hc13f;
aud[3751]=16'hc143;
aud[3752]=16'hc147;
aud[3753]=16'hc14c;
aud[3754]=16'hc150;
aud[3755]=16'hc154;
aud[3756]=16'hc159;
aud[3757]=16'hc15d;
aud[3758]=16'hc162;
aud[3759]=16'hc166;
aud[3760]=16'hc16b;
aud[3761]=16'hc16f;
aud[3762]=16'hc174;
aud[3763]=16'hc178;
aud[3764]=16'hc17d;
aud[3765]=16'hc181;
aud[3766]=16'hc186;
aud[3767]=16'hc18b;
aud[3768]=16'hc18f;
aud[3769]=16'hc194;
aud[3770]=16'hc199;
aud[3771]=16'hc19e;
aud[3772]=16'hc1a2;
aud[3773]=16'hc1a7;
aud[3774]=16'hc1ac;
aud[3775]=16'hc1b1;
aud[3776]=16'hc1b6;
aud[3777]=16'hc1bb;
aud[3778]=16'hc1c0;
aud[3779]=16'hc1c5;
aud[3780]=16'hc1ca;
aud[3781]=16'hc1cf;
aud[3782]=16'hc1d4;
aud[3783]=16'hc1d9;
aud[3784]=16'hc1de;
aud[3785]=16'hc1e3;
aud[3786]=16'hc1e8;
aud[3787]=16'hc1ee;
aud[3788]=16'hc1f3;
aud[3789]=16'hc1f8;
aud[3790]=16'hc1fd;
aud[3791]=16'hc203;
aud[3792]=16'hc208;
aud[3793]=16'hc20d;
aud[3794]=16'hc213;
aud[3795]=16'hc218;
aud[3796]=16'hc21e;
aud[3797]=16'hc223;
aud[3798]=16'hc229;
aud[3799]=16'hc22e;
aud[3800]=16'hc234;
aud[3801]=16'hc239;
aud[3802]=16'hc23f;
aud[3803]=16'hc245;
aud[3804]=16'hc24a;
aud[3805]=16'hc250;
aud[3806]=16'hc256;
aud[3807]=16'hc25c;
aud[3808]=16'hc261;
aud[3809]=16'hc267;
aud[3810]=16'hc26d;
aud[3811]=16'hc273;
aud[3812]=16'hc279;
aud[3813]=16'hc27f;
aud[3814]=16'hc285;
aud[3815]=16'hc28b;
aud[3816]=16'hc291;
aud[3817]=16'hc297;
aud[3818]=16'hc29d;
aud[3819]=16'hc2a3;
aud[3820]=16'hc2a9;
aud[3821]=16'hc2af;
aud[3822]=16'hc2b5;
aud[3823]=16'hc2bb;
aud[3824]=16'hc2c1;
aud[3825]=16'hc2c8;
aud[3826]=16'hc2ce;
aud[3827]=16'hc2d4;
aud[3828]=16'hc2db;
aud[3829]=16'hc2e1;
aud[3830]=16'hc2e7;
aud[3831]=16'hc2ee;
aud[3832]=16'hc2f4;
aud[3833]=16'hc2fb;
aud[3834]=16'hc301;
aud[3835]=16'hc308;
aud[3836]=16'hc30e;
aud[3837]=16'hc315;
aud[3838]=16'hc31b;
aud[3839]=16'hc322;
aud[3840]=16'hc329;
aud[3841]=16'hc32f;
aud[3842]=16'hc336;
aud[3843]=16'hc33d;
aud[3844]=16'hc343;
aud[3845]=16'hc34a;
aud[3846]=16'hc351;
aud[3847]=16'hc358;
aud[3848]=16'hc35f;
aud[3849]=16'hc365;
aud[3850]=16'hc36c;
aud[3851]=16'hc373;
aud[3852]=16'hc37a;
aud[3853]=16'hc381;
aud[3854]=16'hc388;
aud[3855]=16'hc38f;
aud[3856]=16'hc396;
aud[3857]=16'hc39d;
aud[3858]=16'hc3a5;
aud[3859]=16'hc3ac;
aud[3860]=16'hc3b3;
aud[3861]=16'hc3ba;
aud[3862]=16'hc3c1;
aud[3863]=16'hc3c9;
aud[3864]=16'hc3d0;
aud[3865]=16'hc3d7;
aud[3866]=16'hc3df;
aud[3867]=16'hc3e6;
aud[3868]=16'hc3ed;
aud[3869]=16'hc3f5;
aud[3870]=16'hc3fc;
aud[3871]=16'hc404;
aud[3872]=16'hc40b;
aud[3873]=16'hc413;
aud[3874]=16'hc41a;
aud[3875]=16'hc422;
aud[3876]=16'hc429;
aud[3877]=16'hc431;
aud[3878]=16'hc439;
aud[3879]=16'hc440;
aud[3880]=16'hc448;
aud[3881]=16'hc450;
aud[3882]=16'hc457;
aud[3883]=16'hc45f;
aud[3884]=16'hc467;
aud[3885]=16'hc46f;
aud[3886]=16'hc477;
aud[3887]=16'hc47f;
aud[3888]=16'hc486;
aud[3889]=16'hc48e;
aud[3890]=16'hc496;
aud[3891]=16'hc49e;
aud[3892]=16'hc4a6;
aud[3893]=16'hc4ae;
aud[3894]=16'hc4b6;
aud[3895]=16'hc4bf;
aud[3896]=16'hc4c7;
aud[3897]=16'hc4cf;
aud[3898]=16'hc4d7;
aud[3899]=16'hc4df;
aud[3900]=16'hc4e7;
aud[3901]=16'hc4f0;
aud[3902]=16'hc4f8;
aud[3903]=16'hc500;
aud[3904]=16'hc509;
aud[3905]=16'hc511;
aud[3906]=16'hc519;
aud[3907]=16'hc522;
aud[3908]=16'hc52a;
aud[3909]=16'hc533;
aud[3910]=16'hc53b;
aud[3911]=16'hc544;
aud[3912]=16'hc54c;
aud[3913]=16'hc555;
aud[3914]=16'hc55d;
aud[3915]=16'hc566;
aud[3916]=16'hc56e;
aud[3917]=16'hc577;
aud[3918]=16'hc580;
aud[3919]=16'hc588;
aud[3920]=16'hc591;
aud[3921]=16'hc59a;
aud[3922]=16'hc5a3;
aud[3923]=16'hc5ac;
aud[3924]=16'hc5b4;
aud[3925]=16'hc5bd;
aud[3926]=16'hc5c6;
aud[3927]=16'hc5cf;
aud[3928]=16'hc5d8;
aud[3929]=16'hc5e1;
aud[3930]=16'hc5ea;
aud[3931]=16'hc5f3;
aud[3932]=16'hc5fc;
aud[3933]=16'hc605;
aud[3934]=16'hc60e;
aud[3935]=16'hc617;
aud[3936]=16'hc620;
aud[3937]=16'hc62a;
aud[3938]=16'hc633;
aud[3939]=16'hc63c;
aud[3940]=16'hc645;
aud[3941]=16'hc64f;
aud[3942]=16'hc658;
aud[3943]=16'hc661;
aud[3944]=16'hc66b;
aud[3945]=16'hc674;
aud[3946]=16'hc67d;
aud[3947]=16'hc687;
aud[3948]=16'hc690;
aud[3949]=16'hc69a;
aud[3950]=16'hc6a3;
aud[3951]=16'hc6ad;
aud[3952]=16'hc6b6;
aud[3953]=16'hc6c0;
aud[3954]=16'hc6c9;
aud[3955]=16'hc6d3;
aud[3956]=16'hc6dd;
aud[3957]=16'hc6e6;
aud[3958]=16'hc6f0;
aud[3959]=16'hc6fa;
aud[3960]=16'hc703;
aud[3961]=16'hc70d;
aud[3962]=16'hc717;
aud[3963]=16'hc721;
aud[3964]=16'hc72b;
aud[3965]=16'hc735;
aud[3966]=16'hc73f;
aud[3967]=16'hc748;
aud[3968]=16'hc752;
aud[3969]=16'hc75c;
aud[3970]=16'hc766;
aud[3971]=16'hc770;
aud[3972]=16'hc77a;
aud[3973]=16'hc785;
aud[3974]=16'hc78f;
aud[3975]=16'hc799;
aud[3976]=16'hc7a3;
aud[3977]=16'hc7ad;
aud[3978]=16'hc7b7;
aud[3979]=16'hc7c1;
aud[3980]=16'hc7cc;
aud[3981]=16'hc7d6;
aud[3982]=16'hc7e0;
aud[3983]=16'hc7eb;
aud[3984]=16'hc7f5;
aud[3985]=16'hc7ff;
aud[3986]=16'hc80a;
aud[3987]=16'hc814;
aud[3988]=16'hc81f;
aud[3989]=16'hc829;
aud[3990]=16'hc834;
aud[3991]=16'hc83e;
aud[3992]=16'hc849;
aud[3993]=16'hc853;
aud[3994]=16'hc85e;
aud[3995]=16'hc868;
aud[3996]=16'hc873;
aud[3997]=16'hc87e;
aud[3998]=16'hc888;
aud[3999]=16'hc893;
aud[4000]=16'hc89e;
aud[4001]=16'hc8a9;
aud[4002]=16'hc8b3;
aud[4003]=16'hc8be;
aud[4004]=16'hc8c9;
aud[4005]=16'hc8d4;
aud[4006]=16'hc8df;
aud[4007]=16'hc8ea;
aud[4008]=16'hc8f5;
aud[4009]=16'hc8ff;
aud[4010]=16'hc90a;
aud[4011]=16'hc915;
aud[4012]=16'hc920;
aud[4013]=16'hc92c;
aud[4014]=16'hc937;
aud[4015]=16'hc942;
aud[4016]=16'hc94d;
aud[4017]=16'hc958;
aud[4018]=16'hc963;
aud[4019]=16'hc96e;
aud[4020]=16'hc97a;
aud[4021]=16'hc985;
aud[4022]=16'hc990;
aud[4023]=16'hc99b;
aud[4024]=16'hc9a7;
aud[4025]=16'hc9b2;
aud[4026]=16'hc9bd;
aud[4027]=16'hc9c9;
aud[4028]=16'hc9d4;
aud[4029]=16'hc9e0;
aud[4030]=16'hc9eb;
aud[4031]=16'hc9f7;
aud[4032]=16'hca02;
aud[4033]=16'hca0e;
aud[4034]=16'hca19;
aud[4035]=16'hca25;
aud[4036]=16'hca30;
aud[4037]=16'hca3c;
aud[4038]=16'hca48;
aud[4039]=16'hca53;
aud[4040]=16'hca5f;
aud[4041]=16'hca6b;
aud[4042]=16'hca76;
aud[4043]=16'hca82;
aud[4044]=16'hca8e;
aud[4045]=16'hca9a;
aud[4046]=16'hcaa6;
aud[4047]=16'hcab1;
aud[4048]=16'hcabd;
aud[4049]=16'hcac9;
aud[4050]=16'hcad5;
aud[4051]=16'hcae1;
aud[4052]=16'hcaed;
aud[4053]=16'hcaf9;
aud[4054]=16'hcb05;
aud[4055]=16'hcb11;
aud[4056]=16'hcb1d;
aud[4057]=16'hcb29;
aud[4058]=16'hcb35;
aud[4059]=16'hcb42;
aud[4060]=16'hcb4e;
aud[4061]=16'hcb5a;
aud[4062]=16'hcb66;
aud[4063]=16'hcb72;
aud[4064]=16'hcb7f;
aud[4065]=16'hcb8b;
aud[4066]=16'hcb97;
aud[4067]=16'hcba3;
aud[4068]=16'hcbb0;
aud[4069]=16'hcbbc;
aud[4070]=16'hcbc9;
aud[4071]=16'hcbd5;
aud[4072]=16'hcbe1;
aud[4073]=16'hcbee;
aud[4074]=16'hcbfa;
aud[4075]=16'hcc07;
aud[4076]=16'hcc13;
aud[4077]=16'hcc20;
aud[4078]=16'hcc2c;
aud[4079]=16'hcc39;
aud[4080]=16'hcc46;
aud[4081]=16'hcc52;
aud[4082]=16'hcc5f;
aud[4083]=16'hcc6c;
aud[4084]=16'hcc78;
aud[4085]=16'hcc85;
aud[4086]=16'hcc92;
aud[4087]=16'hcc9f;
aud[4088]=16'hccab;
aud[4089]=16'hccb8;
aud[4090]=16'hccc5;
aud[4091]=16'hccd2;
aud[4092]=16'hccdf;
aud[4093]=16'hccec;
aud[4094]=16'hccf9;
aud[4095]=16'hcd06;
aud[4096]=16'hcd13;
aud[4097]=16'hcd20;
aud[4098]=16'hcd2d;
aud[4099]=16'hcd3a;
aud[4100]=16'hcd47;
aud[4101]=16'hcd54;
aud[4102]=16'hcd61;
aud[4103]=16'hcd6e;
aud[4104]=16'hcd7b;
aud[4105]=16'hcd88;
aud[4106]=16'hcd96;
aud[4107]=16'hcda3;
aud[4108]=16'hcdb0;
aud[4109]=16'hcdbd;
aud[4110]=16'hcdcb;
aud[4111]=16'hcdd8;
aud[4112]=16'hcde5;
aud[4113]=16'hcdf3;
aud[4114]=16'hce00;
aud[4115]=16'hce0d;
aud[4116]=16'hce1b;
aud[4117]=16'hce28;
aud[4118]=16'hce36;
aud[4119]=16'hce43;
aud[4120]=16'hce51;
aud[4121]=16'hce5e;
aud[4122]=16'hce6c;
aud[4123]=16'hce79;
aud[4124]=16'hce87;
aud[4125]=16'hce95;
aud[4126]=16'hcea2;
aud[4127]=16'hceb0;
aud[4128]=16'hcebe;
aud[4129]=16'hcecb;
aud[4130]=16'hced9;
aud[4131]=16'hcee7;
aud[4132]=16'hcef5;
aud[4133]=16'hcf02;
aud[4134]=16'hcf10;
aud[4135]=16'hcf1e;
aud[4136]=16'hcf2c;
aud[4137]=16'hcf3a;
aud[4138]=16'hcf48;
aud[4139]=16'hcf56;
aud[4140]=16'hcf63;
aud[4141]=16'hcf71;
aud[4142]=16'hcf7f;
aud[4143]=16'hcf8d;
aud[4144]=16'hcf9b;
aud[4145]=16'hcfa9;
aud[4146]=16'hcfb8;
aud[4147]=16'hcfc6;
aud[4148]=16'hcfd4;
aud[4149]=16'hcfe2;
aud[4150]=16'hcff0;
aud[4151]=16'hcffe;
aud[4152]=16'hd00c;
aud[4153]=16'hd01b;
aud[4154]=16'hd029;
aud[4155]=16'hd037;
aud[4156]=16'hd045;
aud[4157]=16'hd054;
aud[4158]=16'hd062;
aud[4159]=16'hd070;
aud[4160]=16'hd07f;
aud[4161]=16'hd08d;
aud[4162]=16'hd09b;
aud[4163]=16'hd0aa;
aud[4164]=16'hd0b8;
aud[4165]=16'hd0c7;
aud[4166]=16'hd0d5;
aud[4167]=16'hd0e4;
aud[4168]=16'hd0f2;
aud[4169]=16'hd101;
aud[4170]=16'hd10f;
aud[4171]=16'hd11e;
aud[4172]=16'hd12d;
aud[4173]=16'hd13b;
aud[4174]=16'hd14a;
aud[4175]=16'hd159;
aud[4176]=16'hd167;
aud[4177]=16'hd176;
aud[4178]=16'hd185;
aud[4179]=16'hd193;
aud[4180]=16'hd1a2;
aud[4181]=16'hd1b1;
aud[4182]=16'hd1c0;
aud[4183]=16'hd1cf;
aud[4184]=16'hd1de;
aud[4185]=16'hd1ec;
aud[4186]=16'hd1fb;
aud[4187]=16'hd20a;
aud[4188]=16'hd219;
aud[4189]=16'hd228;
aud[4190]=16'hd237;
aud[4191]=16'hd246;
aud[4192]=16'hd255;
aud[4193]=16'hd264;
aud[4194]=16'hd273;
aud[4195]=16'hd282;
aud[4196]=16'hd291;
aud[4197]=16'hd2a0;
aud[4198]=16'hd2b0;
aud[4199]=16'hd2bf;
aud[4200]=16'hd2ce;
aud[4201]=16'hd2dd;
aud[4202]=16'hd2ec;
aud[4203]=16'hd2fc;
aud[4204]=16'hd30b;
aud[4205]=16'hd31a;
aud[4206]=16'hd329;
aud[4207]=16'hd339;
aud[4208]=16'hd348;
aud[4209]=16'hd357;
aud[4210]=16'hd367;
aud[4211]=16'hd376;
aud[4212]=16'hd386;
aud[4213]=16'hd395;
aud[4214]=16'hd3a4;
aud[4215]=16'hd3b4;
aud[4216]=16'hd3c3;
aud[4217]=16'hd3d3;
aud[4218]=16'hd3e2;
aud[4219]=16'hd3f2;
aud[4220]=16'hd402;
aud[4221]=16'hd411;
aud[4222]=16'hd421;
aud[4223]=16'hd430;
aud[4224]=16'hd440;
aud[4225]=16'hd450;
aud[4226]=16'hd45f;
aud[4227]=16'hd46f;
aud[4228]=16'hd47f;
aud[4229]=16'hd48f;
aud[4230]=16'hd49e;
aud[4231]=16'hd4ae;
aud[4232]=16'hd4be;
aud[4233]=16'hd4ce;
aud[4234]=16'hd4de;
aud[4235]=16'hd4ed;
aud[4236]=16'hd4fd;
aud[4237]=16'hd50d;
aud[4238]=16'hd51d;
aud[4239]=16'hd52d;
aud[4240]=16'hd53d;
aud[4241]=16'hd54d;
aud[4242]=16'hd55d;
aud[4243]=16'hd56d;
aud[4244]=16'hd57d;
aud[4245]=16'hd58d;
aud[4246]=16'hd59d;
aud[4247]=16'hd5ad;
aud[4248]=16'hd5bd;
aud[4249]=16'hd5cd;
aud[4250]=16'hd5dd;
aud[4251]=16'hd5ee;
aud[4252]=16'hd5fe;
aud[4253]=16'hd60e;
aud[4254]=16'hd61e;
aud[4255]=16'hd62e;
aud[4256]=16'hd63f;
aud[4257]=16'hd64f;
aud[4258]=16'hd65f;
aud[4259]=16'hd66f;
aud[4260]=16'hd680;
aud[4261]=16'hd690;
aud[4262]=16'hd6a0;
aud[4263]=16'hd6b1;
aud[4264]=16'hd6c1;
aud[4265]=16'hd6d2;
aud[4266]=16'hd6e2;
aud[4267]=16'hd6f2;
aud[4268]=16'hd703;
aud[4269]=16'hd713;
aud[4270]=16'hd724;
aud[4271]=16'hd734;
aud[4272]=16'hd745;
aud[4273]=16'hd756;
aud[4274]=16'hd766;
aud[4275]=16'hd777;
aud[4276]=16'hd787;
aud[4277]=16'hd798;
aud[4278]=16'hd7a9;
aud[4279]=16'hd7b9;
aud[4280]=16'hd7ca;
aud[4281]=16'hd7db;
aud[4282]=16'hd7eb;
aud[4283]=16'hd7fc;
aud[4284]=16'hd80d;
aud[4285]=16'hd81e;
aud[4286]=16'hd82e;
aud[4287]=16'hd83f;
aud[4288]=16'hd850;
aud[4289]=16'hd861;
aud[4290]=16'hd872;
aud[4291]=16'hd882;
aud[4292]=16'hd893;
aud[4293]=16'hd8a4;
aud[4294]=16'hd8b5;
aud[4295]=16'hd8c6;
aud[4296]=16'hd8d7;
aud[4297]=16'hd8e8;
aud[4298]=16'hd8f9;
aud[4299]=16'hd90a;
aud[4300]=16'hd91b;
aud[4301]=16'hd92c;
aud[4302]=16'hd93d;
aud[4303]=16'hd94e;
aud[4304]=16'hd95f;
aud[4305]=16'hd970;
aud[4306]=16'hd982;
aud[4307]=16'hd993;
aud[4308]=16'hd9a4;
aud[4309]=16'hd9b5;
aud[4310]=16'hd9c6;
aud[4311]=16'hd9d7;
aud[4312]=16'hd9e9;
aud[4313]=16'hd9fa;
aud[4314]=16'hda0b;
aud[4315]=16'hda1c;
aud[4316]=16'hda2e;
aud[4317]=16'hda3f;
aud[4318]=16'hda50;
aud[4319]=16'hda62;
aud[4320]=16'hda73;
aud[4321]=16'hda84;
aud[4322]=16'hda96;
aud[4323]=16'hdaa7;
aud[4324]=16'hdab9;
aud[4325]=16'hdaca;
aud[4326]=16'hdadc;
aud[4327]=16'hdaed;
aud[4328]=16'hdaff;
aud[4329]=16'hdb10;
aud[4330]=16'hdb22;
aud[4331]=16'hdb33;
aud[4332]=16'hdb45;
aud[4333]=16'hdb56;
aud[4334]=16'hdb68;
aud[4335]=16'hdb79;
aud[4336]=16'hdb8b;
aud[4337]=16'hdb9d;
aud[4338]=16'hdbae;
aud[4339]=16'hdbc0;
aud[4340]=16'hdbd2;
aud[4341]=16'hdbe3;
aud[4342]=16'hdbf5;
aud[4343]=16'hdc07;
aud[4344]=16'hdc19;
aud[4345]=16'hdc2a;
aud[4346]=16'hdc3c;
aud[4347]=16'hdc4e;
aud[4348]=16'hdc60;
aud[4349]=16'hdc72;
aud[4350]=16'hdc83;
aud[4351]=16'hdc95;
aud[4352]=16'hdca7;
aud[4353]=16'hdcb9;
aud[4354]=16'hdccb;
aud[4355]=16'hdcdd;
aud[4356]=16'hdcef;
aud[4357]=16'hdd01;
aud[4358]=16'hdd13;
aud[4359]=16'hdd25;
aud[4360]=16'hdd37;
aud[4361]=16'hdd49;
aud[4362]=16'hdd5b;
aud[4363]=16'hdd6d;
aud[4364]=16'hdd7f;
aud[4365]=16'hdd91;
aud[4366]=16'hdda3;
aud[4367]=16'hddb5;
aud[4368]=16'hddc7;
aud[4369]=16'hddd9;
aud[4370]=16'hddeb;
aud[4371]=16'hddfe;
aud[4372]=16'hde10;
aud[4373]=16'hde22;
aud[4374]=16'hde34;
aud[4375]=16'hde46;
aud[4376]=16'hde59;
aud[4377]=16'hde6b;
aud[4378]=16'hde7d;
aud[4379]=16'hde8f;
aud[4380]=16'hdea2;
aud[4381]=16'hdeb4;
aud[4382]=16'hdec6;
aud[4383]=16'hded9;
aud[4384]=16'hdeeb;
aud[4385]=16'hdefd;
aud[4386]=16'hdf10;
aud[4387]=16'hdf22;
aud[4388]=16'hdf35;
aud[4389]=16'hdf47;
aud[4390]=16'hdf59;
aud[4391]=16'hdf6c;
aud[4392]=16'hdf7e;
aud[4393]=16'hdf91;
aud[4394]=16'hdfa3;
aud[4395]=16'hdfb6;
aud[4396]=16'hdfc8;
aud[4397]=16'hdfdb;
aud[4398]=16'hdfed;
aud[4399]=16'he000;
aud[4400]=16'he013;
aud[4401]=16'he025;
aud[4402]=16'he038;
aud[4403]=16'he04a;
aud[4404]=16'he05d;
aud[4405]=16'he070;
aud[4406]=16'he082;
aud[4407]=16'he095;
aud[4408]=16'he0a8;
aud[4409]=16'he0ba;
aud[4410]=16'he0cd;
aud[4411]=16'he0e0;
aud[4412]=16'he0f3;
aud[4413]=16'he105;
aud[4414]=16'he118;
aud[4415]=16'he12b;
aud[4416]=16'he13e;
aud[4417]=16'he151;
aud[4418]=16'he163;
aud[4419]=16'he176;
aud[4420]=16'he189;
aud[4421]=16'he19c;
aud[4422]=16'he1af;
aud[4423]=16'he1c2;
aud[4424]=16'he1d5;
aud[4425]=16'he1e8;
aud[4426]=16'he1fa;
aud[4427]=16'he20d;
aud[4428]=16'he220;
aud[4429]=16'he233;
aud[4430]=16'he246;
aud[4431]=16'he259;
aud[4432]=16'he26c;
aud[4433]=16'he27f;
aud[4434]=16'he292;
aud[4435]=16'he2a5;
aud[4436]=16'he2b9;
aud[4437]=16'he2cc;
aud[4438]=16'he2df;
aud[4439]=16'he2f2;
aud[4440]=16'he305;
aud[4441]=16'he318;
aud[4442]=16'he32b;
aud[4443]=16'he33e;
aud[4444]=16'he352;
aud[4445]=16'he365;
aud[4446]=16'he378;
aud[4447]=16'he38b;
aud[4448]=16'he39e;
aud[4449]=16'he3b2;
aud[4450]=16'he3c5;
aud[4451]=16'he3d8;
aud[4452]=16'he3eb;
aud[4453]=16'he3ff;
aud[4454]=16'he412;
aud[4455]=16'he425;
aud[4456]=16'he438;
aud[4457]=16'he44c;
aud[4458]=16'he45f;
aud[4459]=16'he473;
aud[4460]=16'he486;
aud[4461]=16'he499;
aud[4462]=16'he4ad;
aud[4463]=16'he4c0;
aud[4464]=16'he4d3;
aud[4465]=16'he4e7;
aud[4466]=16'he4fa;
aud[4467]=16'he50e;
aud[4468]=16'he521;
aud[4469]=16'he535;
aud[4470]=16'he548;
aud[4471]=16'he55c;
aud[4472]=16'he56f;
aud[4473]=16'he583;
aud[4474]=16'he596;
aud[4475]=16'he5aa;
aud[4476]=16'he5bd;
aud[4477]=16'he5d1;
aud[4478]=16'he5e4;
aud[4479]=16'he5f8;
aud[4480]=16'he60c;
aud[4481]=16'he61f;
aud[4482]=16'he633;
aud[4483]=16'he646;
aud[4484]=16'he65a;
aud[4485]=16'he66e;
aud[4486]=16'he681;
aud[4487]=16'he695;
aud[4488]=16'he6a9;
aud[4489]=16'he6bd;
aud[4490]=16'he6d0;
aud[4491]=16'he6e4;
aud[4492]=16'he6f8;
aud[4493]=16'he70b;
aud[4494]=16'he71f;
aud[4495]=16'he733;
aud[4496]=16'he747;
aud[4497]=16'he75b;
aud[4498]=16'he76e;
aud[4499]=16'he782;
aud[4500]=16'he796;
aud[4501]=16'he7aa;
aud[4502]=16'he7be;
aud[4503]=16'he7d1;
aud[4504]=16'he7e5;
aud[4505]=16'he7f9;
aud[4506]=16'he80d;
aud[4507]=16'he821;
aud[4508]=16'he835;
aud[4509]=16'he849;
aud[4510]=16'he85d;
aud[4511]=16'he871;
aud[4512]=16'he885;
aud[4513]=16'he899;
aud[4514]=16'he8ad;
aud[4515]=16'he8c0;
aud[4516]=16'he8d4;
aud[4517]=16'he8e8;
aud[4518]=16'he8fc;
aud[4519]=16'he910;
aud[4520]=16'he925;
aud[4521]=16'he939;
aud[4522]=16'he94d;
aud[4523]=16'he961;
aud[4524]=16'he975;
aud[4525]=16'he989;
aud[4526]=16'he99d;
aud[4527]=16'he9b1;
aud[4528]=16'he9c5;
aud[4529]=16'he9d9;
aud[4530]=16'he9ed;
aud[4531]=16'hea01;
aud[4532]=16'hea16;
aud[4533]=16'hea2a;
aud[4534]=16'hea3e;
aud[4535]=16'hea52;
aud[4536]=16'hea66;
aud[4537]=16'hea7a;
aud[4538]=16'hea8f;
aud[4539]=16'heaa3;
aud[4540]=16'heab7;
aud[4541]=16'heacb;
aud[4542]=16'heae0;
aud[4543]=16'heaf4;
aud[4544]=16'heb08;
aud[4545]=16'heb1c;
aud[4546]=16'heb31;
aud[4547]=16'heb45;
aud[4548]=16'heb59;
aud[4549]=16'heb6e;
aud[4550]=16'heb82;
aud[4551]=16'heb96;
aud[4552]=16'hebab;
aud[4553]=16'hebbf;
aud[4554]=16'hebd3;
aud[4555]=16'hebe8;
aud[4556]=16'hebfc;
aud[4557]=16'hec10;
aud[4558]=16'hec25;
aud[4559]=16'hec39;
aud[4560]=16'hec4d;
aud[4561]=16'hec62;
aud[4562]=16'hec76;
aud[4563]=16'hec8b;
aud[4564]=16'hec9f;
aud[4565]=16'hecb4;
aud[4566]=16'hecc8;
aud[4567]=16'hecdd;
aud[4568]=16'hecf1;
aud[4569]=16'hed05;
aud[4570]=16'hed1a;
aud[4571]=16'hed2e;
aud[4572]=16'hed43;
aud[4573]=16'hed57;
aud[4574]=16'hed6c;
aud[4575]=16'hed81;
aud[4576]=16'hed95;
aud[4577]=16'hedaa;
aud[4578]=16'hedbe;
aud[4579]=16'hedd3;
aud[4580]=16'hede7;
aud[4581]=16'hedfc;
aud[4582]=16'hee10;
aud[4583]=16'hee25;
aud[4584]=16'hee3a;
aud[4585]=16'hee4e;
aud[4586]=16'hee63;
aud[4587]=16'hee77;
aud[4588]=16'hee8c;
aud[4589]=16'heea1;
aud[4590]=16'heeb5;
aud[4591]=16'heeca;
aud[4592]=16'heedf;
aud[4593]=16'heef3;
aud[4594]=16'hef08;
aud[4595]=16'hef1d;
aud[4596]=16'hef31;
aud[4597]=16'hef46;
aud[4598]=16'hef5b;
aud[4599]=16'hef70;
aud[4600]=16'hef84;
aud[4601]=16'hef99;
aud[4602]=16'hefae;
aud[4603]=16'hefc2;
aud[4604]=16'hefd7;
aud[4605]=16'hefec;
aud[4606]=16'hf001;
aud[4607]=16'hf015;
aud[4608]=16'hf02a;
aud[4609]=16'hf03f;
aud[4610]=16'hf054;
aud[4611]=16'hf069;
aud[4612]=16'hf07d;
aud[4613]=16'hf092;
aud[4614]=16'hf0a7;
aud[4615]=16'hf0bc;
aud[4616]=16'hf0d1;
aud[4617]=16'hf0e6;
aud[4618]=16'hf0fa;
aud[4619]=16'hf10f;
aud[4620]=16'hf124;
aud[4621]=16'hf139;
aud[4622]=16'hf14e;
aud[4623]=16'hf163;
aud[4624]=16'hf178;
aud[4625]=16'hf18c;
aud[4626]=16'hf1a1;
aud[4627]=16'hf1b6;
aud[4628]=16'hf1cb;
aud[4629]=16'hf1e0;
aud[4630]=16'hf1f5;
aud[4631]=16'hf20a;
aud[4632]=16'hf21f;
aud[4633]=16'hf234;
aud[4634]=16'hf249;
aud[4635]=16'hf25e;
aud[4636]=16'hf273;
aud[4637]=16'hf288;
aud[4638]=16'hf29d;
aud[4639]=16'hf2b2;
aud[4640]=16'hf2c7;
aud[4641]=16'hf2dc;
aud[4642]=16'hf2f1;
aud[4643]=16'hf306;
aud[4644]=16'hf31b;
aud[4645]=16'hf330;
aud[4646]=16'hf345;
aud[4647]=16'hf35a;
aud[4648]=16'hf36f;
aud[4649]=16'hf384;
aud[4650]=16'hf399;
aud[4651]=16'hf3ae;
aud[4652]=16'hf3c3;
aud[4653]=16'hf3d8;
aud[4654]=16'hf3ed;
aud[4655]=16'hf402;
aud[4656]=16'hf417;
aud[4657]=16'hf42c;
aud[4658]=16'hf441;
aud[4659]=16'hf456;
aud[4660]=16'hf46b;
aud[4661]=16'hf480;
aud[4662]=16'hf496;
aud[4663]=16'hf4ab;
aud[4664]=16'hf4c0;
aud[4665]=16'hf4d5;
aud[4666]=16'hf4ea;
aud[4667]=16'hf4ff;
aud[4668]=16'hf514;
aud[4669]=16'hf529;
aud[4670]=16'hf53f;
aud[4671]=16'hf554;
aud[4672]=16'hf569;
aud[4673]=16'hf57e;
aud[4674]=16'hf593;
aud[4675]=16'hf5a8;
aud[4676]=16'hf5bd;
aud[4677]=16'hf5d3;
aud[4678]=16'hf5e8;
aud[4679]=16'hf5fd;
aud[4680]=16'hf612;
aud[4681]=16'hf627;
aud[4682]=16'hf63d;
aud[4683]=16'hf652;
aud[4684]=16'hf667;
aud[4685]=16'hf67c;
aud[4686]=16'hf691;
aud[4687]=16'hf6a7;
aud[4688]=16'hf6bc;
aud[4689]=16'hf6d1;
aud[4690]=16'hf6e6;
aud[4691]=16'hf6fb;
aud[4692]=16'hf711;
aud[4693]=16'hf726;
aud[4694]=16'hf73b;
aud[4695]=16'hf750;
aud[4696]=16'hf766;
aud[4697]=16'hf77b;
aud[4698]=16'hf790;
aud[4699]=16'hf7a5;
aud[4700]=16'hf7bb;
aud[4701]=16'hf7d0;
aud[4702]=16'hf7e5;
aud[4703]=16'hf7fb;
aud[4704]=16'hf810;
aud[4705]=16'hf825;
aud[4706]=16'hf83a;
aud[4707]=16'hf850;
aud[4708]=16'hf865;
aud[4709]=16'hf87a;
aud[4710]=16'hf890;
aud[4711]=16'hf8a5;
aud[4712]=16'hf8ba;
aud[4713]=16'hf8cf;
aud[4714]=16'hf8e5;
aud[4715]=16'hf8fa;
aud[4716]=16'hf90f;
aud[4717]=16'hf925;
aud[4718]=16'hf93a;
aud[4719]=16'hf94f;
aud[4720]=16'hf965;
aud[4721]=16'hf97a;
aud[4722]=16'hf98f;
aud[4723]=16'hf9a5;
aud[4724]=16'hf9ba;
aud[4725]=16'hf9cf;
aud[4726]=16'hf9e5;
aud[4727]=16'hf9fa;
aud[4728]=16'hfa0f;
aud[4729]=16'hfa25;
aud[4730]=16'hfa3a;
aud[4731]=16'hfa50;
aud[4732]=16'hfa65;
aud[4733]=16'hfa7a;
aud[4734]=16'hfa90;
aud[4735]=16'hfaa5;
aud[4736]=16'hfaba;
aud[4737]=16'hfad0;
aud[4738]=16'hfae5;
aud[4739]=16'hfafb;
aud[4740]=16'hfb10;
aud[4741]=16'hfb25;
aud[4742]=16'hfb3b;
aud[4743]=16'hfb50;
aud[4744]=16'hfb65;
aud[4745]=16'hfb7b;
aud[4746]=16'hfb90;
aud[4747]=16'hfba6;
aud[4748]=16'hfbbb;
aud[4749]=16'hfbd0;
aud[4750]=16'hfbe6;
aud[4751]=16'hfbfb;
aud[4752]=16'hfc11;
aud[4753]=16'hfc26;
aud[4754]=16'hfc3b;
aud[4755]=16'hfc51;
aud[4756]=16'hfc66;
aud[4757]=16'hfc7c;
aud[4758]=16'hfc91;
aud[4759]=16'hfca7;
aud[4760]=16'hfcbc;
aud[4761]=16'hfcd1;
aud[4762]=16'hfce7;
aud[4763]=16'hfcfc;
aud[4764]=16'hfd12;
aud[4765]=16'hfd27;
aud[4766]=16'hfd3c;
aud[4767]=16'hfd52;
aud[4768]=16'hfd67;
aud[4769]=16'hfd7d;
aud[4770]=16'hfd92;
aud[4771]=16'hfda8;
aud[4772]=16'hfdbd;
aud[4773]=16'hfdd2;
aud[4774]=16'hfde8;
aud[4775]=16'hfdfd;
aud[4776]=16'hfe13;
aud[4777]=16'hfe28;
aud[4778]=16'hfe3e;
aud[4779]=16'hfe53;
aud[4780]=16'hfe69;
aud[4781]=16'hfe7e;
aud[4782]=16'hfe93;
aud[4783]=16'hfea9;
aud[4784]=16'hfebe;
aud[4785]=16'hfed4;
aud[4786]=16'hfee9;
aud[4787]=16'hfeff;
aud[4788]=16'hff14;
aud[4789]=16'hff2a;
aud[4790]=16'hff3f;
aud[4791]=16'hff54;
aud[4792]=16'hff6a;
aud[4793]=16'hff7f;
aud[4794]=16'hff95;
aud[4795]=16'hffaa;
aud[4796]=16'hffc0;
aud[4797]=16'hffd5;
aud[4798]=16'hffeb;
aud[4799]=16'h0;
aud[4800]=16'h15;
aud[4801]=16'h2b;
aud[4802]=16'h40;
aud[4803]=16'h56;
aud[4804]=16'h6b;
aud[4805]=16'h81;
aud[4806]=16'h96;
aud[4807]=16'hac;
aud[4808]=16'hc1;
aud[4809]=16'hd6;
aud[4810]=16'hec;
aud[4811]=16'h101;
aud[4812]=16'h117;
aud[4813]=16'h12c;
aud[4814]=16'h142;
aud[4815]=16'h157;
aud[4816]=16'h16d;
aud[4817]=16'h182;
aud[4818]=16'h197;
aud[4819]=16'h1ad;
aud[4820]=16'h1c2;
aud[4821]=16'h1d8;
aud[4822]=16'h1ed;
aud[4823]=16'h203;
aud[4824]=16'h218;
aud[4825]=16'h22e;
aud[4826]=16'h243;
aud[4827]=16'h258;
aud[4828]=16'h26e;
aud[4829]=16'h283;
aud[4830]=16'h299;
aud[4831]=16'h2ae;
aud[4832]=16'h2c4;
aud[4833]=16'h2d9;
aud[4834]=16'h2ee;
aud[4835]=16'h304;
aud[4836]=16'h319;
aud[4837]=16'h32f;
aud[4838]=16'h344;
aud[4839]=16'h359;
aud[4840]=16'h36f;
aud[4841]=16'h384;
aud[4842]=16'h39a;
aud[4843]=16'h3af;
aud[4844]=16'h3c5;
aud[4845]=16'h3da;
aud[4846]=16'h3ef;
aud[4847]=16'h405;
aud[4848]=16'h41a;
aud[4849]=16'h430;
aud[4850]=16'h445;
aud[4851]=16'h45a;
aud[4852]=16'h470;
aud[4853]=16'h485;
aud[4854]=16'h49b;
aud[4855]=16'h4b0;
aud[4856]=16'h4c5;
aud[4857]=16'h4db;
aud[4858]=16'h4f0;
aud[4859]=16'h505;
aud[4860]=16'h51b;
aud[4861]=16'h530;
aud[4862]=16'h546;
aud[4863]=16'h55b;
aud[4864]=16'h570;
aud[4865]=16'h586;
aud[4866]=16'h59b;
aud[4867]=16'h5b0;
aud[4868]=16'h5c6;
aud[4869]=16'h5db;
aud[4870]=16'h5f1;
aud[4871]=16'h606;
aud[4872]=16'h61b;
aud[4873]=16'h631;
aud[4874]=16'h646;
aud[4875]=16'h65b;
aud[4876]=16'h671;
aud[4877]=16'h686;
aud[4878]=16'h69b;
aud[4879]=16'h6b1;
aud[4880]=16'h6c6;
aud[4881]=16'h6db;
aud[4882]=16'h6f1;
aud[4883]=16'h706;
aud[4884]=16'h71b;
aud[4885]=16'h731;
aud[4886]=16'h746;
aud[4887]=16'h75b;
aud[4888]=16'h770;
aud[4889]=16'h786;
aud[4890]=16'h79b;
aud[4891]=16'h7b0;
aud[4892]=16'h7c6;
aud[4893]=16'h7db;
aud[4894]=16'h7f0;
aud[4895]=16'h805;
aud[4896]=16'h81b;
aud[4897]=16'h830;
aud[4898]=16'h845;
aud[4899]=16'h85b;
aud[4900]=16'h870;
aud[4901]=16'h885;
aud[4902]=16'h89a;
aud[4903]=16'h8b0;
aud[4904]=16'h8c5;
aud[4905]=16'h8da;
aud[4906]=16'h8ef;
aud[4907]=16'h905;
aud[4908]=16'h91a;
aud[4909]=16'h92f;
aud[4910]=16'h944;
aud[4911]=16'h959;
aud[4912]=16'h96f;
aud[4913]=16'h984;
aud[4914]=16'h999;
aud[4915]=16'h9ae;
aud[4916]=16'h9c3;
aud[4917]=16'h9d9;
aud[4918]=16'h9ee;
aud[4919]=16'ha03;
aud[4920]=16'ha18;
aud[4921]=16'ha2d;
aud[4922]=16'ha43;
aud[4923]=16'ha58;
aud[4924]=16'ha6d;
aud[4925]=16'ha82;
aud[4926]=16'ha97;
aud[4927]=16'haac;
aud[4928]=16'hac1;
aud[4929]=16'had7;
aud[4930]=16'haec;
aud[4931]=16'hb01;
aud[4932]=16'hb16;
aud[4933]=16'hb2b;
aud[4934]=16'hb40;
aud[4935]=16'hb55;
aud[4936]=16'hb6a;
aud[4937]=16'hb80;
aud[4938]=16'hb95;
aud[4939]=16'hbaa;
aud[4940]=16'hbbf;
aud[4941]=16'hbd4;
aud[4942]=16'hbe9;
aud[4943]=16'hbfe;
aud[4944]=16'hc13;
aud[4945]=16'hc28;
aud[4946]=16'hc3d;
aud[4947]=16'hc52;
aud[4948]=16'hc67;
aud[4949]=16'hc7c;
aud[4950]=16'hc91;
aud[4951]=16'hca6;
aud[4952]=16'hcbb;
aud[4953]=16'hcd0;
aud[4954]=16'hce5;
aud[4955]=16'hcfa;
aud[4956]=16'hd0f;
aud[4957]=16'hd24;
aud[4958]=16'hd39;
aud[4959]=16'hd4e;
aud[4960]=16'hd63;
aud[4961]=16'hd78;
aud[4962]=16'hd8d;
aud[4963]=16'hda2;
aud[4964]=16'hdb7;
aud[4965]=16'hdcc;
aud[4966]=16'hde1;
aud[4967]=16'hdf6;
aud[4968]=16'he0b;
aud[4969]=16'he20;
aud[4970]=16'he35;
aud[4971]=16'he4a;
aud[4972]=16'he5f;
aud[4973]=16'he74;
aud[4974]=16'he88;
aud[4975]=16'he9d;
aud[4976]=16'heb2;
aud[4977]=16'hec7;
aud[4978]=16'hedc;
aud[4979]=16'hef1;
aud[4980]=16'hf06;
aud[4981]=16'hf1a;
aud[4982]=16'hf2f;
aud[4983]=16'hf44;
aud[4984]=16'hf59;
aud[4985]=16'hf6e;
aud[4986]=16'hf83;
aud[4987]=16'hf97;
aud[4988]=16'hfac;
aud[4989]=16'hfc1;
aud[4990]=16'hfd6;
aud[4991]=16'hfeb;
aud[4992]=16'hfff;
aud[4993]=16'h1014;
aud[4994]=16'h1029;
aud[4995]=16'h103e;
aud[4996]=16'h1052;
aud[4997]=16'h1067;
aud[4998]=16'h107c;
aud[4999]=16'h1090;
aud[5000]=16'h10a5;
aud[5001]=16'h10ba;
aud[5002]=16'h10cf;
aud[5003]=16'h10e3;
aud[5004]=16'h10f8;
aud[5005]=16'h110d;
aud[5006]=16'h1121;
aud[5007]=16'h1136;
aud[5008]=16'h114b;
aud[5009]=16'h115f;
aud[5010]=16'h1174;
aud[5011]=16'h1189;
aud[5012]=16'h119d;
aud[5013]=16'h11b2;
aud[5014]=16'h11c6;
aud[5015]=16'h11db;
aud[5016]=16'h11f0;
aud[5017]=16'h1204;
aud[5018]=16'h1219;
aud[5019]=16'h122d;
aud[5020]=16'h1242;
aud[5021]=16'h1256;
aud[5022]=16'h126b;
aud[5023]=16'h127f;
aud[5024]=16'h1294;
aud[5025]=16'h12a9;
aud[5026]=16'h12bd;
aud[5027]=16'h12d2;
aud[5028]=16'h12e6;
aud[5029]=16'h12fb;
aud[5030]=16'h130f;
aud[5031]=16'h1323;
aud[5032]=16'h1338;
aud[5033]=16'h134c;
aud[5034]=16'h1361;
aud[5035]=16'h1375;
aud[5036]=16'h138a;
aud[5037]=16'h139e;
aud[5038]=16'h13b3;
aud[5039]=16'h13c7;
aud[5040]=16'h13db;
aud[5041]=16'h13f0;
aud[5042]=16'h1404;
aud[5043]=16'h1418;
aud[5044]=16'h142d;
aud[5045]=16'h1441;
aud[5046]=16'h1455;
aud[5047]=16'h146a;
aud[5048]=16'h147e;
aud[5049]=16'h1492;
aud[5050]=16'h14a7;
aud[5051]=16'h14bb;
aud[5052]=16'h14cf;
aud[5053]=16'h14e4;
aud[5054]=16'h14f8;
aud[5055]=16'h150c;
aud[5056]=16'h1520;
aud[5057]=16'h1535;
aud[5058]=16'h1549;
aud[5059]=16'h155d;
aud[5060]=16'h1571;
aud[5061]=16'h1586;
aud[5062]=16'h159a;
aud[5063]=16'h15ae;
aud[5064]=16'h15c2;
aud[5065]=16'h15d6;
aud[5066]=16'h15ea;
aud[5067]=16'h15ff;
aud[5068]=16'h1613;
aud[5069]=16'h1627;
aud[5070]=16'h163b;
aud[5071]=16'h164f;
aud[5072]=16'h1663;
aud[5073]=16'h1677;
aud[5074]=16'h168b;
aud[5075]=16'h169f;
aud[5076]=16'h16b3;
aud[5077]=16'h16c7;
aud[5078]=16'h16db;
aud[5079]=16'h16f0;
aud[5080]=16'h1704;
aud[5081]=16'h1718;
aud[5082]=16'h172c;
aud[5083]=16'h1740;
aud[5084]=16'h1753;
aud[5085]=16'h1767;
aud[5086]=16'h177b;
aud[5087]=16'h178f;
aud[5088]=16'h17a3;
aud[5089]=16'h17b7;
aud[5090]=16'h17cb;
aud[5091]=16'h17df;
aud[5092]=16'h17f3;
aud[5093]=16'h1807;
aud[5094]=16'h181b;
aud[5095]=16'h182f;
aud[5096]=16'h1842;
aud[5097]=16'h1856;
aud[5098]=16'h186a;
aud[5099]=16'h187e;
aud[5100]=16'h1892;
aud[5101]=16'h18a5;
aud[5102]=16'h18b9;
aud[5103]=16'h18cd;
aud[5104]=16'h18e1;
aud[5105]=16'h18f5;
aud[5106]=16'h1908;
aud[5107]=16'h191c;
aud[5108]=16'h1930;
aud[5109]=16'h1943;
aud[5110]=16'h1957;
aud[5111]=16'h196b;
aud[5112]=16'h197f;
aud[5113]=16'h1992;
aud[5114]=16'h19a6;
aud[5115]=16'h19ba;
aud[5116]=16'h19cd;
aud[5117]=16'h19e1;
aud[5118]=16'h19f4;
aud[5119]=16'h1a08;
aud[5120]=16'h1a1c;
aud[5121]=16'h1a2f;
aud[5122]=16'h1a43;
aud[5123]=16'h1a56;
aud[5124]=16'h1a6a;
aud[5125]=16'h1a7d;
aud[5126]=16'h1a91;
aud[5127]=16'h1aa4;
aud[5128]=16'h1ab8;
aud[5129]=16'h1acb;
aud[5130]=16'h1adf;
aud[5131]=16'h1af2;
aud[5132]=16'h1b06;
aud[5133]=16'h1b19;
aud[5134]=16'h1b2d;
aud[5135]=16'h1b40;
aud[5136]=16'h1b53;
aud[5137]=16'h1b67;
aud[5138]=16'h1b7a;
aud[5139]=16'h1b8d;
aud[5140]=16'h1ba1;
aud[5141]=16'h1bb4;
aud[5142]=16'h1bc8;
aud[5143]=16'h1bdb;
aud[5144]=16'h1bee;
aud[5145]=16'h1c01;
aud[5146]=16'h1c15;
aud[5147]=16'h1c28;
aud[5148]=16'h1c3b;
aud[5149]=16'h1c4e;
aud[5150]=16'h1c62;
aud[5151]=16'h1c75;
aud[5152]=16'h1c88;
aud[5153]=16'h1c9b;
aud[5154]=16'h1cae;
aud[5155]=16'h1cc2;
aud[5156]=16'h1cd5;
aud[5157]=16'h1ce8;
aud[5158]=16'h1cfb;
aud[5159]=16'h1d0e;
aud[5160]=16'h1d21;
aud[5161]=16'h1d34;
aud[5162]=16'h1d47;
aud[5163]=16'h1d5b;
aud[5164]=16'h1d6e;
aud[5165]=16'h1d81;
aud[5166]=16'h1d94;
aud[5167]=16'h1da7;
aud[5168]=16'h1dba;
aud[5169]=16'h1dcd;
aud[5170]=16'h1de0;
aud[5171]=16'h1df3;
aud[5172]=16'h1e06;
aud[5173]=16'h1e18;
aud[5174]=16'h1e2b;
aud[5175]=16'h1e3e;
aud[5176]=16'h1e51;
aud[5177]=16'h1e64;
aud[5178]=16'h1e77;
aud[5179]=16'h1e8a;
aud[5180]=16'h1e9d;
aud[5181]=16'h1eaf;
aud[5182]=16'h1ec2;
aud[5183]=16'h1ed5;
aud[5184]=16'h1ee8;
aud[5185]=16'h1efb;
aud[5186]=16'h1f0d;
aud[5187]=16'h1f20;
aud[5188]=16'h1f33;
aud[5189]=16'h1f46;
aud[5190]=16'h1f58;
aud[5191]=16'h1f6b;
aud[5192]=16'h1f7e;
aud[5193]=16'h1f90;
aud[5194]=16'h1fa3;
aud[5195]=16'h1fb6;
aud[5196]=16'h1fc8;
aud[5197]=16'h1fdb;
aud[5198]=16'h1fed;
aud[5199]=16'h2000;
aud[5200]=16'h2013;
aud[5201]=16'h2025;
aud[5202]=16'h2038;
aud[5203]=16'h204a;
aud[5204]=16'h205d;
aud[5205]=16'h206f;
aud[5206]=16'h2082;
aud[5207]=16'h2094;
aud[5208]=16'h20a7;
aud[5209]=16'h20b9;
aud[5210]=16'h20cb;
aud[5211]=16'h20de;
aud[5212]=16'h20f0;
aud[5213]=16'h2103;
aud[5214]=16'h2115;
aud[5215]=16'h2127;
aud[5216]=16'h213a;
aud[5217]=16'h214c;
aud[5218]=16'h215e;
aud[5219]=16'h2171;
aud[5220]=16'h2183;
aud[5221]=16'h2195;
aud[5222]=16'h21a7;
aud[5223]=16'h21ba;
aud[5224]=16'h21cc;
aud[5225]=16'h21de;
aud[5226]=16'h21f0;
aud[5227]=16'h2202;
aud[5228]=16'h2215;
aud[5229]=16'h2227;
aud[5230]=16'h2239;
aud[5231]=16'h224b;
aud[5232]=16'h225d;
aud[5233]=16'h226f;
aud[5234]=16'h2281;
aud[5235]=16'h2293;
aud[5236]=16'h22a5;
aud[5237]=16'h22b7;
aud[5238]=16'h22c9;
aud[5239]=16'h22db;
aud[5240]=16'h22ed;
aud[5241]=16'h22ff;
aud[5242]=16'h2311;
aud[5243]=16'h2323;
aud[5244]=16'h2335;
aud[5245]=16'h2347;
aud[5246]=16'h2359;
aud[5247]=16'h236b;
aud[5248]=16'h237d;
aud[5249]=16'h238e;
aud[5250]=16'h23a0;
aud[5251]=16'h23b2;
aud[5252]=16'h23c4;
aud[5253]=16'h23d6;
aud[5254]=16'h23e7;
aud[5255]=16'h23f9;
aud[5256]=16'h240b;
aud[5257]=16'h241d;
aud[5258]=16'h242e;
aud[5259]=16'h2440;
aud[5260]=16'h2452;
aud[5261]=16'h2463;
aud[5262]=16'h2475;
aud[5263]=16'h2487;
aud[5264]=16'h2498;
aud[5265]=16'h24aa;
aud[5266]=16'h24bb;
aud[5267]=16'h24cd;
aud[5268]=16'h24de;
aud[5269]=16'h24f0;
aud[5270]=16'h2501;
aud[5271]=16'h2513;
aud[5272]=16'h2524;
aud[5273]=16'h2536;
aud[5274]=16'h2547;
aud[5275]=16'h2559;
aud[5276]=16'h256a;
aud[5277]=16'h257c;
aud[5278]=16'h258d;
aud[5279]=16'h259e;
aud[5280]=16'h25b0;
aud[5281]=16'h25c1;
aud[5282]=16'h25d2;
aud[5283]=16'h25e4;
aud[5284]=16'h25f5;
aud[5285]=16'h2606;
aud[5286]=16'h2617;
aud[5287]=16'h2629;
aud[5288]=16'h263a;
aud[5289]=16'h264b;
aud[5290]=16'h265c;
aud[5291]=16'h266d;
aud[5292]=16'h267e;
aud[5293]=16'h2690;
aud[5294]=16'h26a1;
aud[5295]=16'h26b2;
aud[5296]=16'h26c3;
aud[5297]=16'h26d4;
aud[5298]=16'h26e5;
aud[5299]=16'h26f6;
aud[5300]=16'h2707;
aud[5301]=16'h2718;
aud[5302]=16'h2729;
aud[5303]=16'h273a;
aud[5304]=16'h274b;
aud[5305]=16'h275c;
aud[5306]=16'h276d;
aud[5307]=16'h277e;
aud[5308]=16'h278e;
aud[5309]=16'h279f;
aud[5310]=16'h27b0;
aud[5311]=16'h27c1;
aud[5312]=16'h27d2;
aud[5313]=16'h27e2;
aud[5314]=16'h27f3;
aud[5315]=16'h2804;
aud[5316]=16'h2815;
aud[5317]=16'h2825;
aud[5318]=16'h2836;
aud[5319]=16'h2847;
aud[5320]=16'h2857;
aud[5321]=16'h2868;
aud[5322]=16'h2879;
aud[5323]=16'h2889;
aud[5324]=16'h289a;
aud[5325]=16'h28aa;
aud[5326]=16'h28bb;
aud[5327]=16'h28cc;
aud[5328]=16'h28dc;
aud[5329]=16'h28ed;
aud[5330]=16'h28fd;
aud[5331]=16'h290e;
aud[5332]=16'h291e;
aud[5333]=16'h292e;
aud[5334]=16'h293f;
aud[5335]=16'h294f;
aud[5336]=16'h2960;
aud[5337]=16'h2970;
aud[5338]=16'h2980;
aud[5339]=16'h2991;
aud[5340]=16'h29a1;
aud[5341]=16'h29b1;
aud[5342]=16'h29c1;
aud[5343]=16'h29d2;
aud[5344]=16'h29e2;
aud[5345]=16'h29f2;
aud[5346]=16'h2a02;
aud[5347]=16'h2a12;
aud[5348]=16'h2a23;
aud[5349]=16'h2a33;
aud[5350]=16'h2a43;
aud[5351]=16'h2a53;
aud[5352]=16'h2a63;
aud[5353]=16'h2a73;
aud[5354]=16'h2a83;
aud[5355]=16'h2a93;
aud[5356]=16'h2aa3;
aud[5357]=16'h2ab3;
aud[5358]=16'h2ac3;
aud[5359]=16'h2ad3;
aud[5360]=16'h2ae3;
aud[5361]=16'h2af3;
aud[5362]=16'h2b03;
aud[5363]=16'h2b13;
aud[5364]=16'h2b22;
aud[5365]=16'h2b32;
aud[5366]=16'h2b42;
aud[5367]=16'h2b52;
aud[5368]=16'h2b62;
aud[5369]=16'h2b71;
aud[5370]=16'h2b81;
aud[5371]=16'h2b91;
aud[5372]=16'h2ba1;
aud[5373]=16'h2bb0;
aud[5374]=16'h2bc0;
aud[5375]=16'h2bd0;
aud[5376]=16'h2bdf;
aud[5377]=16'h2bef;
aud[5378]=16'h2bfe;
aud[5379]=16'h2c0e;
aud[5380]=16'h2c1e;
aud[5381]=16'h2c2d;
aud[5382]=16'h2c3d;
aud[5383]=16'h2c4c;
aud[5384]=16'h2c5c;
aud[5385]=16'h2c6b;
aud[5386]=16'h2c7a;
aud[5387]=16'h2c8a;
aud[5388]=16'h2c99;
aud[5389]=16'h2ca9;
aud[5390]=16'h2cb8;
aud[5391]=16'h2cc7;
aud[5392]=16'h2cd7;
aud[5393]=16'h2ce6;
aud[5394]=16'h2cf5;
aud[5395]=16'h2d04;
aud[5396]=16'h2d14;
aud[5397]=16'h2d23;
aud[5398]=16'h2d32;
aud[5399]=16'h2d41;
aud[5400]=16'h2d50;
aud[5401]=16'h2d60;
aud[5402]=16'h2d6f;
aud[5403]=16'h2d7e;
aud[5404]=16'h2d8d;
aud[5405]=16'h2d9c;
aud[5406]=16'h2dab;
aud[5407]=16'h2dba;
aud[5408]=16'h2dc9;
aud[5409]=16'h2dd8;
aud[5410]=16'h2de7;
aud[5411]=16'h2df6;
aud[5412]=16'h2e05;
aud[5413]=16'h2e14;
aud[5414]=16'h2e22;
aud[5415]=16'h2e31;
aud[5416]=16'h2e40;
aud[5417]=16'h2e4f;
aud[5418]=16'h2e5e;
aud[5419]=16'h2e6d;
aud[5420]=16'h2e7b;
aud[5421]=16'h2e8a;
aud[5422]=16'h2e99;
aud[5423]=16'h2ea7;
aud[5424]=16'h2eb6;
aud[5425]=16'h2ec5;
aud[5426]=16'h2ed3;
aud[5427]=16'h2ee2;
aud[5428]=16'h2ef1;
aud[5429]=16'h2eff;
aud[5430]=16'h2f0e;
aud[5431]=16'h2f1c;
aud[5432]=16'h2f2b;
aud[5433]=16'h2f39;
aud[5434]=16'h2f48;
aud[5435]=16'h2f56;
aud[5436]=16'h2f65;
aud[5437]=16'h2f73;
aud[5438]=16'h2f81;
aud[5439]=16'h2f90;
aud[5440]=16'h2f9e;
aud[5441]=16'h2fac;
aud[5442]=16'h2fbb;
aud[5443]=16'h2fc9;
aud[5444]=16'h2fd7;
aud[5445]=16'h2fe5;
aud[5446]=16'h2ff4;
aud[5447]=16'h3002;
aud[5448]=16'h3010;
aud[5449]=16'h301e;
aud[5450]=16'h302c;
aud[5451]=16'h303a;
aud[5452]=16'h3048;
aud[5453]=16'h3057;
aud[5454]=16'h3065;
aud[5455]=16'h3073;
aud[5456]=16'h3081;
aud[5457]=16'h308f;
aud[5458]=16'h309d;
aud[5459]=16'h30aa;
aud[5460]=16'h30b8;
aud[5461]=16'h30c6;
aud[5462]=16'h30d4;
aud[5463]=16'h30e2;
aud[5464]=16'h30f0;
aud[5465]=16'h30fe;
aud[5466]=16'h310b;
aud[5467]=16'h3119;
aud[5468]=16'h3127;
aud[5469]=16'h3135;
aud[5470]=16'h3142;
aud[5471]=16'h3150;
aud[5472]=16'h315e;
aud[5473]=16'h316b;
aud[5474]=16'h3179;
aud[5475]=16'h3187;
aud[5476]=16'h3194;
aud[5477]=16'h31a2;
aud[5478]=16'h31af;
aud[5479]=16'h31bd;
aud[5480]=16'h31ca;
aud[5481]=16'h31d8;
aud[5482]=16'h31e5;
aud[5483]=16'h31f3;
aud[5484]=16'h3200;
aud[5485]=16'h320d;
aud[5486]=16'h321b;
aud[5487]=16'h3228;
aud[5488]=16'h3235;
aud[5489]=16'h3243;
aud[5490]=16'h3250;
aud[5491]=16'h325d;
aud[5492]=16'h326a;
aud[5493]=16'h3278;
aud[5494]=16'h3285;
aud[5495]=16'h3292;
aud[5496]=16'h329f;
aud[5497]=16'h32ac;
aud[5498]=16'h32b9;
aud[5499]=16'h32c6;
aud[5500]=16'h32d3;
aud[5501]=16'h32e0;
aud[5502]=16'h32ed;
aud[5503]=16'h32fa;
aud[5504]=16'h3307;
aud[5505]=16'h3314;
aud[5506]=16'h3321;
aud[5507]=16'h332e;
aud[5508]=16'h333b;
aud[5509]=16'h3348;
aud[5510]=16'h3355;
aud[5511]=16'h3361;
aud[5512]=16'h336e;
aud[5513]=16'h337b;
aud[5514]=16'h3388;
aud[5515]=16'h3394;
aud[5516]=16'h33a1;
aud[5517]=16'h33ae;
aud[5518]=16'h33ba;
aud[5519]=16'h33c7;
aud[5520]=16'h33d4;
aud[5521]=16'h33e0;
aud[5522]=16'h33ed;
aud[5523]=16'h33f9;
aud[5524]=16'h3406;
aud[5525]=16'h3412;
aud[5526]=16'h341f;
aud[5527]=16'h342b;
aud[5528]=16'h3437;
aud[5529]=16'h3444;
aud[5530]=16'h3450;
aud[5531]=16'h345d;
aud[5532]=16'h3469;
aud[5533]=16'h3475;
aud[5534]=16'h3481;
aud[5535]=16'h348e;
aud[5536]=16'h349a;
aud[5537]=16'h34a6;
aud[5538]=16'h34b2;
aud[5539]=16'h34be;
aud[5540]=16'h34cb;
aud[5541]=16'h34d7;
aud[5542]=16'h34e3;
aud[5543]=16'h34ef;
aud[5544]=16'h34fb;
aud[5545]=16'h3507;
aud[5546]=16'h3513;
aud[5547]=16'h351f;
aud[5548]=16'h352b;
aud[5549]=16'h3537;
aud[5550]=16'h3543;
aud[5551]=16'h354f;
aud[5552]=16'h355a;
aud[5553]=16'h3566;
aud[5554]=16'h3572;
aud[5555]=16'h357e;
aud[5556]=16'h358a;
aud[5557]=16'h3595;
aud[5558]=16'h35a1;
aud[5559]=16'h35ad;
aud[5560]=16'h35b8;
aud[5561]=16'h35c4;
aud[5562]=16'h35d0;
aud[5563]=16'h35db;
aud[5564]=16'h35e7;
aud[5565]=16'h35f2;
aud[5566]=16'h35fe;
aud[5567]=16'h3609;
aud[5568]=16'h3615;
aud[5569]=16'h3620;
aud[5570]=16'h362c;
aud[5571]=16'h3637;
aud[5572]=16'h3643;
aud[5573]=16'h364e;
aud[5574]=16'h3659;
aud[5575]=16'h3665;
aud[5576]=16'h3670;
aud[5577]=16'h367b;
aud[5578]=16'h3686;
aud[5579]=16'h3692;
aud[5580]=16'h369d;
aud[5581]=16'h36a8;
aud[5582]=16'h36b3;
aud[5583]=16'h36be;
aud[5584]=16'h36c9;
aud[5585]=16'h36d4;
aud[5586]=16'h36e0;
aud[5587]=16'h36eb;
aud[5588]=16'h36f6;
aud[5589]=16'h3701;
aud[5590]=16'h370b;
aud[5591]=16'h3716;
aud[5592]=16'h3721;
aud[5593]=16'h372c;
aud[5594]=16'h3737;
aud[5595]=16'h3742;
aud[5596]=16'h374d;
aud[5597]=16'h3757;
aud[5598]=16'h3762;
aud[5599]=16'h376d;
aud[5600]=16'h3778;
aud[5601]=16'h3782;
aud[5602]=16'h378d;
aud[5603]=16'h3798;
aud[5604]=16'h37a2;
aud[5605]=16'h37ad;
aud[5606]=16'h37b7;
aud[5607]=16'h37c2;
aud[5608]=16'h37cc;
aud[5609]=16'h37d7;
aud[5610]=16'h37e1;
aud[5611]=16'h37ec;
aud[5612]=16'h37f6;
aud[5613]=16'h3801;
aud[5614]=16'h380b;
aud[5615]=16'h3815;
aud[5616]=16'h3820;
aud[5617]=16'h382a;
aud[5618]=16'h3834;
aud[5619]=16'h383f;
aud[5620]=16'h3849;
aud[5621]=16'h3853;
aud[5622]=16'h385d;
aud[5623]=16'h3867;
aud[5624]=16'h3871;
aud[5625]=16'h387b;
aud[5626]=16'h3886;
aud[5627]=16'h3890;
aud[5628]=16'h389a;
aud[5629]=16'h38a4;
aud[5630]=16'h38ae;
aud[5631]=16'h38b8;
aud[5632]=16'h38c1;
aud[5633]=16'h38cb;
aud[5634]=16'h38d5;
aud[5635]=16'h38df;
aud[5636]=16'h38e9;
aud[5637]=16'h38f3;
aud[5638]=16'h38fd;
aud[5639]=16'h3906;
aud[5640]=16'h3910;
aud[5641]=16'h391a;
aud[5642]=16'h3923;
aud[5643]=16'h392d;
aud[5644]=16'h3937;
aud[5645]=16'h3940;
aud[5646]=16'h394a;
aud[5647]=16'h3953;
aud[5648]=16'h395d;
aud[5649]=16'h3966;
aud[5650]=16'h3970;
aud[5651]=16'h3979;
aud[5652]=16'h3983;
aud[5653]=16'h398c;
aud[5654]=16'h3995;
aud[5655]=16'h399f;
aud[5656]=16'h39a8;
aud[5657]=16'h39b1;
aud[5658]=16'h39bb;
aud[5659]=16'h39c4;
aud[5660]=16'h39cd;
aud[5661]=16'h39d6;
aud[5662]=16'h39e0;
aud[5663]=16'h39e9;
aud[5664]=16'h39f2;
aud[5665]=16'h39fb;
aud[5666]=16'h3a04;
aud[5667]=16'h3a0d;
aud[5668]=16'h3a16;
aud[5669]=16'h3a1f;
aud[5670]=16'h3a28;
aud[5671]=16'h3a31;
aud[5672]=16'h3a3a;
aud[5673]=16'h3a43;
aud[5674]=16'h3a4c;
aud[5675]=16'h3a54;
aud[5676]=16'h3a5d;
aud[5677]=16'h3a66;
aud[5678]=16'h3a6f;
aud[5679]=16'h3a78;
aud[5680]=16'h3a80;
aud[5681]=16'h3a89;
aud[5682]=16'h3a92;
aud[5683]=16'h3a9a;
aud[5684]=16'h3aa3;
aud[5685]=16'h3aab;
aud[5686]=16'h3ab4;
aud[5687]=16'h3abc;
aud[5688]=16'h3ac5;
aud[5689]=16'h3acd;
aud[5690]=16'h3ad6;
aud[5691]=16'h3ade;
aud[5692]=16'h3ae7;
aud[5693]=16'h3aef;
aud[5694]=16'h3af7;
aud[5695]=16'h3b00;
aud[5696]=16'h3b08;
aud[5697]=16'h3b10;
aud[5698]=16'h3b19;
aud[5699]=16'h3b21;
aud[5700]=16'h3b29;
aud[5701]=16'h3b31;
aud[5702]=16'h3b39;
aud[5703]=16'h3b41;
aud[5704]=16'h3b4a;
aud[5705]=16'h3b52;
aud[5706]=16'h3b5a;
aud[5707]=16'h3b62;
aud[5708]=16'h3b6a;
aud[5709]=16'h3b72;
aud[5710]=16'h3b7a;
aud[5711]=16'h3b81;
aud[5712]=16'h3b89;
aud[5713]=16'h3b91;
aud[5714]=16'h3b99;
aud[5715]=16'h3ba1;
aud[5716]=16'h3ba9;
aud[5717]=16'h3bb0;
aud[5718]=16'h3bb8;
aud[5719]=16'h3bc0;
aud[5720]=16'h3bc7;
aud[5721]=16'h3bcf;
aud[5722]=16'h3bd7;
aud[5723]=16'h3bde;
aud[5724]=16'h3be6;
aud[5725]=16'h3bed;
aud[5726]=16'h3bf5;
aud[5727]=16'h3bfc;
aud[5728]=16'h3c04;
aud[5729]=16'h3c0b;
aud[5730]=16'h3c13;
aud[5731]=16'h3c1a;
aud[5732]=16'h3c21;
aud[5733]=16'h3c29;
aud[5734]=16'h3c30;
aud[5735]=16'h3c37;
aud[5736]=16'h3c3f;
aud[5737]=16'h3c46;
aud[5738]=16'h3c4d;
aud[5739]=16'h3c54;
aud[5740]=16'h3c5b;
aud[5741]=16'h3c63;
aud[5742]=16'h3c6a;
aud[5743]=16'h3c71;
aud[5744]=16'h3c78;
aud[5745]=16'h3c7f;
aud[5746]=16'h3c86;
aud[5747]=16'h3c8d;
aud[5748]=16'h3c94;
aud[5749]=16'h3c9b;
aud[5750]=16'h3ca1;
aud[5751]=16'h3ca8;
aud[5752]=16'h3caf;
aud[5753]=16'h3cb6;
aud[5754]=16'h3cbd;
aud[5755]=16'h3cc3;
aud[5756]=16'h3cca;
aud[5757]=16'h3cd1;
aud[5758]=16'h3cd7;
aud[5759]=16'h3cde;
aud[5760]=16'h3ce5;
aud[5761]=16'h3ceb;
aud[5762]=16'h3cf2;
aud[5763]=16'h3cf8;
aud[5764]=16'h3cff;
aud[5765]=16'h3d05;
aud[5766]=16'h3d0c;
aud[5767]=16'h3d12;
aud[5768]=16'h3d19;
aud[5769]=16'h3d1f;
aud[5770]=16'h3d25;
aud[5771]=16'h3d2c;
aud[5772]=16'h3d32;
aud[5773]=16'h3d38;
aud[5774]=16'h3d3f;
aud[5775]=16'h3d45;
aud[5776]=16'h3d4b;
aud[5777]=16'h3d51;
aud[5778]=16'h3d57;
aud[5779]=16'h3d5d;
aud[5780]=16'h3d63;
aud[5781]=16'h3d69;
aud[5782]=16'h3d6f;
aud[5783]=16'h3d75;
aud[5784]=16'h3d7b;
aud[5785]=16'h3d81;
aud[5786]=16'h3d87;
aud[5787]=16'h3d8d;
aud[5788]=16'h3d93;
aud[5789]=16'h3d99;
aud[5790]=16'h3d9f;
aud[5791]=16'h3da4;
aud[5792]=16'h3daa;
aud[5793]=16'h3db0;
aud[5794]=16'h3db6;
aud[5795]=16'h3dbb;
aud[5796]=16'h3dc1;
aud[5797]=16'h3dc7;
aud[5798]=16'h3dcc;
aud[5799]=16'h3dd2;
aud[5800]=16'h3dd7;
aud[5801]=16'h3ddd;
aud[5802]=16'h3de2;
aud[5803]=16'h3de8;
aud[5804]=16'h3ded;
aud[5805]=16'h3df3;
aud[5806]=16'h3df8;
aud[5807]=16'h3dfd;
aud[5808]=16'h3e03;
aud[5809]=16'h3e08;
aud[5810]=16'h3e0d;
aud[5811]=16'h3e12;
aud[5812]=16'h3e18;
aud[5813]=16'h3e1d;
aud[5814]=16'h3e22;
aud[5815]=16'h3e27;
aud[5816]=16'h3e2c;
aud[5817]=16'h3e31;
aud[5818]=16'h3e36;
aud[5819]=16'h3e3b;
aud[5820]=16'h3e40;
aud[5821]=16'h3e45;
aud[5822]=16'h3e4a;
aud[5823]=16'h3e4f;
aud[5824]=16'h3e54;
aud[5825]=16'h3e59;
aud[5826]=16'h3e5e;
aud[5827]=16'h3e62;
aud[5828]=16'h3e67;
aud[5829]=16'h3e6c;
aud[5830]=16'h3e71;
aud[5831]=16'h3e75;
aud[5832]=16'h3e7a;
aud[5833]=16'h3e7f;
aud[5834]=16'h3e83;
aud[5835]=16'h3e88;
aud[5836]=16'h3e8c;
aud[5837]=16'h3e91;
aud[5838]=16'h3e95;
aud[5839]=16'h3e9a;
aud[5840]=16'h3e9e;
aud[5841]=16'h3ea3;
aud[5842]=16'h3ea7;
aud[5843]=16'h3eac;
aud[5844]=16'h3eb0;
aud[5845]=16'h3eb4;
aud[5846]=16'h3eb9;
aud[5847]=16'h3ebd;
aud[5848]=16'h3ec1;
aud[5849]=16'h3ec5;
aud[5850]=16'h3ec9;
aud[5851]=16'h3ecd;
aud[5852]=16'h3ed2;
aud[5853]=16'h3ed6;
aud[5854]=16'h3eda;
aud[5855]=16'h3ede;
aud[5856]=16'h3ee2;
aud[5857]=16'h3ee6;
aud[5858]=16'h3eea;
aud[5859]=16'h3eee;
aud[5860]=16'h3ef2;
aud[5861]=16'h3ef5;
aud[5862]=16'h3ef9;
aud[5863]=16'h3efd;
aud[5864]=16'h3f01;
aud[5865]=16'h3f05;
aud[5866]=16'h3f08;
aud[5867]=16'h3f0c;
aud[5868]=16'h3f10;
aud[5869]=16'h3f13;
aud[5870]=16'h3f17;
aud[5871]=16'h3f1b;
aud[5872]=16'h3f1e;
aud[5873]=16'h3f22;
aud[5874]=16'h3f25;
aud[5875]=16'h3f29;
aud[5876]=16'h3f2c;
aud[5877]=16'h3f30;
aud[5878]=16'h3f33;
aud[5879]=16'h3f36;
aud[5880]=16'h3f3a;
aud[5881]=16'h3f3d;
aud[5882]=16'h3f40;
aud[5883]=16'h3f43;
aud[5884]=16'h3f47;
aud[5885]=16'h3f4a;
aud[5886]=16'h3f4d;
aud[5887]=16'h3f50;
aud[5888]=16'h3f53;
aud[5889]=16'h3f56;
aud[5890]=16'h3f5a;
aud[5891]=16'h3f5d;
aud[5892]=16'h3f60;
aud[5893]=16'h3f63;
aud[5894]=16'h3f65;
aud[5895]=16'h3f68;
aud[5896]=16'h3f6b;
aud[5897]=16'h3f6e;
aud[5898]=16'h3f71;
aud[5899]=16'h3f74;
aud[5900]=16'h3f77;
aud[5901]=16'h3f79;
aud[5902]=16'h3f7c;
aud[5903]=16'h3f7f;
aud[5904]=16'h3f81;
aud[5905]=16'h3f84;
aud[5906]=16'h3f87;
aud[5907]=16'h3f89;
aud[5908]=16'h3f8c;
aud[5909]=16'h3f8e;
aud[5910]=16'h3f91;
aud[5911]=16'h3f93;
aud[5912]=16'h3f96;
aud[5913]=16'h3f98;
aud[5914]=16'h3f9b;
aud[5915]=16'h3f9d;
aud[5916]=16'h3f9f;
aud[5917]=16'h3fa2;
aud[5918]=16'h3fa4;
aud[5919]=16'h3fa6;
aud[5920]=16'h3fa8;
aud[5921]=16'h3fab;
aud[5922]=16'h3fad;
aud[5923]=16'h3faf;
aud[5924]=16'h3fb1;
aud[5925]=16'h3fb3;
aud[5926]=16'h3fb5;
aud[5927]=16'h3fb7;
aud[5928]=16'h3fb9;
aud[5929]=16'h3fbb;
aud[5930]=16'h3fbd;
aud[5931]=16'h3fbf;
aud[5932]=16'h3fc1;
aud[5933]=16'h3fc3;
aud[5934]=16'h3fc5;
aud[5935]=16'h3fc7;
aud[5936]=16'h3fc8;
aud[5937]=16'h3fca;
aud[5938]=16'h3fcc;
aud[5939]=16'h3fcd;
aud[5940]=16'h3fcf;
aud[5941]=16'h3fd1;
aud[5942]=16'h3fd2;
aud[5943]=16'h3fd4;
aud[5944]=16'h3fd6;
aud[5945]=16'h3fd7;
aud[5946]=16'h3fd9;
aud[5947]=16'h3fda;
aud[5948]=16'h3fdc;
aud[5949]=16'h3fdd;
aud[5950]=16'h3fde;
aud[5951]=16'h3fe0;
aud[5952]=16'h3fe1;
aud[5953]=16'h3fe2;
aud[5954]=16'h3fe4;
aud[5955]=16'h3fe5;
aud[5956]=16'h3fe6;
aud[5957]=16'h3fe7;
aud[5958]=16'h3fe8;
aud[5959]=16'h3fea;
aud[5960]=16'h3feb;
aud[5961]=16'h3fec;
aud[5962]=16'h3fed;
aud[5963]=16'h3fee;
aud[5964]=16'h3fef;
aud[5965]=16'h3ff0;
aud[5966]=16'h3ff1;
aud[5967]=16'h3ff2;
aud[5968]=16'h3ff3;
aud[5969]=16'h3ff3;
aud[5970]=16'h3ff4;
aud[5971]=16'h3ff5;
aud[5972]=16'h3ff6;
aud[5973]=16'h3ff7;
aud[5974]=16'h3ff7;
aud[5975]=16'h3ff8;
aud[5976]=16'h3ff9;
aud[5977]=16'h3ff9;
aud[5978]=16'h3ffa;
aud[5979]=16'h3ffa;
aud[5980]=16'h3ffb;
aud[5981]=16'h3ffb;
aud[5982]=16'h3ffc;
aud[5983]=16'h3ffc;
aud[5984]=16'h3ffd;
aud[5985]=16'h3ffd;
aud[5986]=16'h3ffe;
aud[5987]=16'h3ffe;
aud[5988]=16'h3ffe;
aud[5989]=16'h3fff;
aud[5990]=16'h3fff;
aud[5991]=16'h3fff;
aud[5992]=16'h3fff;
aud[5993]=16'h3fff;
aud[5994]=16'h4000;
aud[5995]=16'h4000;
aud[5996]=16'h4000;
aud[5997]=16'h4000;
aud[5998]=16'h4000;
aud[5999]=16'h4000;
aud[6000]=16'h4000;
aud[6001]=16'h4000;
aud[6002]=16'h4000;
aud[6003]=16'h4000;
aud[6004]=16'h4000;
aud[6005]=16'h3fff;
aud[6006]=16'h3fff;
aud[6007]=16'h3fff;
aud[6008]=16'h3fff;
aud[6009]=16'h3fff;
aud[6010]=16'h3ffe;
aud[6011]=16'h3ffe;
aud[6012]=16'h3ffe;
aud[6013]=16'h3ffd;
aud[6014]=16'h3ffd;
aud[6015]=16'h3ffc;
aud[6016]=16'h3ffc;
aud[6017]=16'h3ffb;
aud[6018]=16'h3ffb;
aud[6019]=16'h3ffa;
aud[6020]=16'h3ffa;
aud[6021]=16'h3ff9;
aud[6022]=16'h3ff9;
aud[6023]=16'h3ff8;
aud[6024]=16'h3ff7;
aud[6025]=16'h3ff7;
aud[6026]=16'h3ff6;
aud[6027]=16'h3ff5;
aud[6028]=16'h3ff4;
aud[6029]=16'h3ff3;
aud[6030]=16'h3ff3;
aud[6031]=16'h3ff2;
aud[6032]=16'h3ff1;
aud[6033]=16'h3ff0;
aud[6034]=16'h3fef;
aud[6035]=16'h3fee;
aud[6036]=16'h3fed;
aud[6037]=16'h3fec;
aud[6038]=16'h3feb;
aud[6039]=16'h3fea;
aud[6040]=16'h3fe8;
aud[6041]=16'h3fe7;
aud[6042]=16'h3fe6;
aud[6043]=16'h3fe5;
aud[6044]=16'h3fe4;
aud[6045]=16'h3fe2;
aud[6046]=16'h3fe1;
aud[6047]=16'h3fe0;
aud[6048]=16'h3fde;
aud[6049]=16'h3fdd;
aud[6050]=16'h3fdc;
aud[6051]=16'h3fda;
aud[6052]=16'h3fd9;
aud[6053]=16'h3fd7;
aud[6054]=16'h3fd6;
aud[6055]=16'h3fd4;
aud[6056]=16'h3fd2;
aud[6057]=16'h3fd1;
aud[6058]=16'h3fcf;
aud[6059]=16'h3fcd;
aud[6060]=16'h3fcc;
aud[6061]=16'h3fca;
aud[6062]=16'h3fc8;
aud[6063]=16'h3fc7;
aud[6064]=16'h3fc5;
aud[6065]=16'h3fc3;
aud[6066]=16'h3fc1;
aud[6067]=16'h3fbf;
aud[6068]=16'h3fbd;
aud[6069]=16'h3fbb;
aud[6070]=16'h3fb9;
aud[6071]=16'h3fb7;
aud[6072]=16'h3fb5;
aud[6073]=16'h3fb3;
aud[6074]=16'h3fb1;
aud[6075]=16'h3faf;
aud[6076]=16'h3fad;
aud[6077]=16'h3fab;
aud[6078]=16'h3fa8;
aud[6079]=16'h3fa6;
aud[6080]=16'h3fa4;
aud[6081]=16'h3fa2;
aud[6082]=16'h3f9f;
aud[6083]=16'h3f9d;
aud[6084]=16'h3f9b;
aud[6085]=16'h3f98;
aud[6086]=16'h3f96;
aud[6087]=16'h3f93;
aud[6088]=16'h3f91;
aud[6089]=16'h3f8e;
aud[6090]=16'h3f8c;
aud[6091]=16'h3f89;
aud[6092]=16'h3f87;
aud[6093]=16'h3f84;
aud[6094]=16'h3f81;
aud[6095]=16'h3f7f;
aud[6096]=16'h3f7c;
aud[6097]=16'h3f79;
aud[6098]=16'h3f77;
aud[6099]=16'h3f74;
aud[6100]=16'h3f71;
aud[6101]=16'h3f6e;
aud[6102]=16'h3f6b;
aud[6103]=16'h3f68;
aud[6104]=16'h3f65;
aud[6105]=16'h3f63;
aud[6106]=16'h3f60;
aud[6107]=16'h3f5d;
aud[6108]=16'h3f5a;
aud[6109]=16'h3f56;
aud[6110]=16'h3f53;
aud[6111]=16'h3f50;
aud[6112]=16'h3f4d;
aud[6113]=16'h3f4a;
aud[6114]=16'h3f47;
aud[6115]=16'h3f43;
aud[6116]=16'h3f40;
aud[6117]=16'h3f3d;
aud[6118]=16'h3f3a;
aud[6119]=16'h3f36;
aud[6120]=16'h3f33;
aud[6121]=16'h3f30;
aud[6122]=16'h3f2c;
aud[6123]=16'h3f29;
aud[6124]=16'h3f25;
aud[6125]=16'h3f22;
aud[6126]=16'h3f1e;
aud[6127]=16'h3f1b;
aud[6128]=16'h3f17;
aud[6129]=16'h3f13;
aud[6130]=16'h3f10;
aud[6131]=16'h3f0c;
aud[6132]=16'h3f08;
aud[6133]=16'h3f05;
aud[6134]=16'h3f01;
aud[6135]=16'h3efd;
aud[6136]=16'h3ef9;
aud[6137]=16'h3ef5;
aud[6138]=16'h3ef2;
aud[6139]=16'h3eee;
aud[6140]=16'h3eea;
aud[6141]=16'h3ee6;
aud[6142]=16'h3ee2;
aud[6143]=16'h3ede;
aud[6144]=16'h3eda;
aud[6145]=16'h3ed6;
aud[6146]=16'h3ed2;
aud[6147]=16'h3ecd;
aud[6148]=16'h3ec9;
aud[6149]=16'h3ec5;
aud[6150]=16'h3ec1;
aud[6151]=16'h3ebd;
aud[6152]=16'h3eb9;
aud[6153]=16'h3eb4;
aud[6154]=16'h3eb0;
aud[6155]=16'h3eac;
aud[6156]=16'h3ea7;
aud[6157]=16'h3ea3;
aud[6158]=16'h3e9e;
aud[6159]=16'h3e9a;
aud[6160]=16'h3e95;
aud[6161]=16'h3e91;
aud[6162]=16'h3e8c;
aud[6163]=16'h3e88;
aud[6164]=16'h3e83;
aud[6165]=16'h3e7f;
aud[6166]=16'h3e7a;
aud[6167]=16'h3e75;
aud[6168]=16'h3e71;
aud[6169]=16'h3e6c;
aud[6170]=16'h3e67;
aud[6171]=16'h3e62;
aud[6172]=16'h3e5e;
aud[6173]=16'h3e59;
aud[6174]=16'h3e54;
aud[6175]=16'h3e4f;
aud[6176]=16'h3e4a;
aud[6177]=16'h3e45;
aud[6178]=16'h3e40;
aud[6179]=16'h3e3b;
aud[6180]=16'h3e36;
aud[6181]=16'h3e31;
aud[6182]=16'h3e2c;
aud[6183]=16'h3e27;
aud[6184]=16'h3e22;
aud[6185]=16'h3e1d;
aud[6186]=16'h3e18;
aud[6187]=16'h3e12;
aud[6188]=16'h3e0d;
aud[6189]=16'h3e08;
aud[6190]=16'h3e03;
aud[6191]=16'h3dfd;
aud[6192]=16'h3df8;
aud[6193]=16'h3df3;
aud[6194]=16'h3ded;
aud[6195]=16'h3de8;
aud[6196]=16'h3de2;
aud[6197]=16'h3ddd;
aud[6198]=16'h3dd7;
aud[6199]=16'h3dd2;
aud[6200]=16'h3dcc;
aud[6201]=16'h3dc7;
aud[6202]=16'h3dc1;
aud[6203]=16'h3dbb;
aud[6204]=16'h3db6;
aud[6205]=16'h3db0;
aud[6206]=16'h3daa;
aud[6207]=16'h3da4;
aud[6208]=16'h3d9f;
aud[6209]=16'h3d99;
aud[6210]=16'h3d93;
aud[6211]=16'h3d8d;
aud[6212]=16'h3d87;
aud[6213]=16'h3d81;
aud[6214]=16'h3d7b;
aud[6215]=16'h3d75;
aud[6216]=16'h3d6f;
aud[6217]=16'h3d69;
aud[6218]=16'h3d63;
aud[6219]=16'h3d5d;
aud[6220]=16'h3d57;
aud[6221]=16'h3d51;
aud[6222]=16'h3d4b;
aud[6223]=16'h3d45;
aud[6224]=16'h3d3f;
aud[6225]=16'h3d38;
aud[6226]=16'h3d32;
aud[6227]=16'h3d2c;
aud[6228]=16'h3d25;
aud[6229]=16'h3d1f;
aud[6230]=16'h3d19;
aud[6231]=16'h3d12;
aud[6232]=16'h3d0c;
aud[6233]=16'h3d05;
aud[6234]=16'h3cff;
aud[6235]=16'h3cf8;
aud[6236]=16'h3cf2;
aud[6237]=16'h3ceb;
aud[6238]=16'h3ce5;
aud[6239]=16'h3cde;
aud[6240]=16'h3cd7;
aud[6241]=16'h3cd1;
aud[6242]=16'h3cca;
aud[6243]=16'h3cc3;
aud[6244]=16'h3cbd;
aud[6245]=16'h3cb6;
aud[6246]=16'h3caf;
aud[6247]=16'h3ca8;
aud[6248]=16'h3ca1;
aud[6249]=16'h3c9b;
aud[6250]=16'h3c94;
aud[6251]=16'h3c8d;
aud[6252]=16'h3c86;
aud[6253]=16'h3c7f;
aud[6254]=16'h3c78;
aud[6255]=16'h3c71;
aud[6256]=16'h3c6a;
aud[6257]=16'h3c63;
aud[6258]=16'h3c5b;
aud[6259]=16'h3c54;
aud[6260]=16'h3c4d;
aud[6261]=16'h3c46;
aud[6262]=16'h3c3f;
aud[6263]=16'h3c37;
aud[6264]=16'h3c30;
aud[6265]=16'h3c29;
aud[6266]=16'h3c21;
aud[6267]=16'h3c1a;
aud[6268]=16'h3c13;
aud[6269]=16'h3c0b;
aud[6270]=16'h3c04;
aud[6271]=16'h3bfc;
aud[6272]=16'h3bf5;
aud[6273]=16'h3bed;
aud[6274]=16'h3be6;
aud[6275]=16'h3bde;
aud[6276]=16'h3bd7;
aud[6277]=16'h3bcf;
aud[6278]=16'h3bc7;
aud[6279]=16'h3bc0;
aud[6280]=16'h3bb8;
aud[6281]=16'h3bb0;
aud[6282]=16'h3ba9;
aud[6283]=16'h3ba1;
aud[6284]=16'h3b99;
aud[6285]=16'h3b91;
aud[6286]=16'h3b89;
aud[6287]=16'h3b81;
aud[6288]=16'h3b7a;
aud[6289]=16'h3b72;
aud[6290]=16'h3b6a;
aud[6291]=16'h3b62;
aud[6292]=16'h3b5a;
aud[6293]=16'h3b52;
aud[6294]=16'h3b4a;
aud[6295]=16'h3b41;
aud[6296]=16'h3b39;
aud[6297]=16'h3b31;
aud[6298]=16'h3b29;
aud[6299]=16'h3b21;
aud[6300]=16'h3b19;
aud[6301]=16'h3b10;
aud[6302]=16'h3b08;
aud[6303]=16'h3b00;
aud[6304]=16'h3af7;
aud[6305]=16'h3aef;
aud[6306]=16'h3ae7;
aud[6307]=16'h3ade;
aud[6308]=16'h3ad6;
aud[6309]=16'h3acd;
aud[6310]=16'h3ac5;
aud[6311]=16'h3abc;
aud[6312]=16'h3ab4;
aud[6313]=16'h3aab;
aud[6314]=16'h3aa3;
aud[6315]=16'h3a9a;
aud[6316]=16'h3a92;
aud[6317]=16'h3a89;
aud[6318]=16'h3a80;
aud[6319]=16'h3a78;
aud[6320]=16'h3a6f;
aud[6321]=16'h3a66;
aud[6322]=16'h3a5d;
aud[6323]=16'h3a54;
aud[6324]=16'h3a4c;
aud[6325]=16'h3a43;
aud[6326]=16'h3a3a;
aud[6327]=16'h3a31;
aud[6328]=16'h3a28;
aud[6329]=16'h3a1f;
aud[6330]=16'h3a16;
aud[6331]=16'h3a0d;
aud[6332]=16'h3a04;
aud[6333]=16'h39fb;
aud[6334]=16'h39f2;
aud[6335]=16'h39e9;
aud[6336]=16'h39e0;
aud[6337]=16'h39d6;
aud[6338]=16'h39cd;
aud[6339]=16'h39c4;
aud[6340]=16'h39bb;
aud[6341]=16'h39b1;
aud[6342]=16'h39a8;
aud[6343]=16'h399f;
aud[6344]=16'h3995;
aud[6345]=16'h398c;
aud[6346]=16'h3983;
aud[6347]=16'h3979;
aud[6348]=16'h3970;
aud[6349]=16'h3966;
aud[6350]=16'h395d;
aud[6351]=16'h3953;
aud[6352]=16'h394a;
aud[6353]=16'h3940;
aud[6354]=16'h3937;
aud[6355]=16'h392d;
aud[6356]=16'h3923;
aud[6357]=16'h391a;
aud[6358]=16'h3910;
aud[6359]=16'h3906;
aud[6360]=16'h38fd;
aud[6361]=16'h38f3;
aud[6362]=16'h38e9;
aud[6363]=16'h38df;
aud[6364]=16'h38d5;
aud[6365]=16'h38cb;
aud[6366]=16'h38c1;
aud[6367]=16'h38b8;
aud[6368]=16'h38ae;
aud[6369]=16'h38a4;
aud[6370]=16'h389a;
aud[6371]=16'h3890;
aud[6372]=16'h3886;
aud[6373]=16'h387b;
aud[6374]=16'h3871;
aud[6375]=16'h3867;
aud[6376]=16'h385d;
aud[6377]=16'h3853;
aud[6378]=16'h3849;
aud[6379]=16'h383f;
aud[6380]=16'h3834;
aud[6381]=16'h382a;
aud[6382]=16'h3820;
aud[6383]=16'h3815;
aud[6384]=16'h380b;
aud[6385]=16'h3801;
aud[6386]=16'h37f6;
aud[6387]=16'h37ec;
aud[6388]=16'h37e1;
aud[6389]=16'h37d7;
aud[6390]=16'h37cc;
aud[6391]=16'h37c2;
aud[6392]=16'h37b7;
aud[6393]=16'h37ad;
aud[6394]=16'h37a2;
aud[6395]=16'h3798;
aud[6396]=16'h378d;
aud[6397]=16'h3782;
aud[6398]=16'h3778;
aud[6399]=16'h376d;
aud[6400]=16'h3762;
aud[6401]=16'h3757;
aud[6402]=16'h374d;
aud[6403]=16'h3742;
aud[6404]=16'h3737;
aud[6405]=16'h372c;
aud[6406]=16'h3721;
aud[6407]=16'h3716;
aud[6408]=16'h370b;
aud[6409]=16'h3701;
aud[6410]=16'h36f6;
aud[6411]=16'h36eb;
aud[6412]=16'h36e0;
aud[6413]=16'h36d4;
aud[6414]=16'h36c9;
aud[6415]=16'h36be;
aud[6416]=16'h36b3;
aud[6417]=16'h36a8;
aud[6418]=16'h369d;
aud[6419]=16'h3692;
aud[6420]=16'h3686;
aud[6421]=16'h367b;
aud[6422]=16'h3670;
aud[6423]=16'h3665;
aud[6424]=16'h3659;
aud[6425]=16'h364e;
aud[6426]=16'h3643;
aud[6427]=16'h3637;
aud[6428]=16'h362c;
aud[6429]=16'h3620;
aud[6430]=16'h3615;
aud[6431]=16'h3609;
aud[6432]=16'h35fe;
aud[6433]=16'h35f2;
aud[6434]=16'h35e7;
aud[6435]=16'h35db;
aud[6436]=16'h35d0;
aud[6437]=16'h35c4;
aud[6438]=16'h35b8;
aud[6439]=16'h35ad;
aud[6440]=16'h35a1;
aud[6441]=16'h3595;
aud[6442]=16'h358a;
aud[6443]=16'h357e;
aud[6444]=16'h3572;
aud[6445]=16'h3566;
aud[6446]=16'h355a;
aud[6447]=16'h354f;
aud[6448]=16'h3543;
aud[6449]=16'h3537;
aud[6450]=16'h352b;
aud[6451]=16'h351f;
aud[6452]=16'h3513;
aud[6453]=16'h3507;
aud[6454]=16'h34fb;
aud[6455]=16'h34ef;
aud[6456]=16'h34e3;
aud[6457]=16'h34d7;
aud[6458]=16'h34cb;
aud[6459]=16'h34be;
aud[6460]=16'h34b2;
aud[6461]=16'h34a6;
aud[6462]=16'h349a;
aud[6463]=16'h348e;
aud[6464]=16'h3481;
aud[6465]=16'h3475;
aud[6466]=16'h3469;
aud[6467]=16'h345d;
aud[6468]=16'h3450;
aud[6469]=16'h3444;
aud[6470]=16'h3437;
aud[6471]=16'h342b;
aud[6472]=16'h341f;
aud[6473]=16'h3412;
aud[6474]=16'h3406;
aud[6475]=16'h33f9;
aud[6476]=16'h33ed;
aud[6477]=16'h33e0;
aud[6478]=16'h33d4;
aud[6479]=16'h33c7;
aud[6480]=16'h33ba;
aud[6481]=16'h33ae;
aud[6482]=16'h33a1;
aud[6483]=16'h3394;
aud[6484]=16'h3388;
aud[6485]=16'h337b;
aud[6486]=16'h336e;
aud[6487]=16'h3361;
aud[6488]=16'h3355;
aud[6489]=16'h3348;
aud[6490]=16'h333b;
aud[6491]=16'h332e;
aud[6492]=16'h3321;
aud[6493]=16'h3314;
aud[6494]=16'h3307;
aud[6495]=16'h32fa;
aud[6496]=16'h32ed;
aud[6497]=16'h32e0;
aud[6498]=16'h32d3;
aud[6499]=16'h32c6;
aud[6500]=16'h32b9;
aud[6501]=16'h32ac;
aud[6502]=16'h329f;
aud[6503]=16'h3292;
aud[6504]=16'h3285;
aud[6505]=16'h3278;
aud[6506]=16'h326a;
aud[6507]=16'h325d;
aud[6508]=16'h3250;
aud[6509]=16'h3243;
aud[6510]=16'h3235;
aud[6511]=16'h3228;
aud[6512]=16'h321b;
aud[6513]=16'h320d;
aud[6514]=16'h3200;
aud[6515]=16'h31f3;
aud[6516]=16'h31e5;
aud[6517]=16'h31d8;
aud[6518]=16'h31ca;
aud[6519]=16'h31bd;
aud[6520]=16'h31af;
aud[6521]=16'h31a2;
aud[6522]=16'h3194;
aud[6523]=16'h3187;
aud[6524]=16'h3179;
aud[6525]=16'h316b;
aud[6526]=16'h315e;
aud[6527]=16'h3150;
aud[6528]=16'h3142;
aud[6529]=16'h3135;
aud[6530]=16'h3127;
aud[6531]=16'h3119;
aud[6532]=16'h310b;
aud[6533]=16'h30fe;
aud[6534]=16'h30f0;
aud[6535]=16'h30e2;
aud[6536]=16'h30d4;
aud[6537]=16'h30c6;
aud[6538]=16'h30b8;
aud[6539]=16'h30aa;
aud[6540]=16'h309d;
aud[6541]=16'h308f;
aud[6542]=16'h3081;
aud[6543]=16'h3073;
aud[6544]=16'h3065;
aud[6545]=16'h3057;
aud[6546]=16'h3048;
aud[6547]=16'h303a;
aud[6548]=16'h302c;
aud[6549]=16'h301e;
aud[6550]=16'h3010;
aud[6551]=16'h3002;
aud[6552]=16'h2ff4;
aud[6553]=16'h2fe5;
aud[6554]=16'h2fd7;
aud[6555]=16'h2fc9;
aud[6556]=16'h2fbb;
aud[6557]=16'h2fac;
aud[6558]=16'h2f9e;
aud[6559]=16'h2f90;
aud[6560]=16'h2f81;
aud[6561]=16'h2f73;
aud[6562]=16'h2f65;
aud[6563]=16'h2f56;
aud[6564]=16'h2f48;
aud[6565]=16'h2f39;
aud[6566]=16'h2f2b;
aud[6567]=16'h2f1c;
aud[6568]=16'h2f0e;
aud[6569]=16'h2eff;
aud[6570]=16'h2ef1;
aud[6571]=16'h2ee2;
aud[6572]=16'h2ed3;
aud[6573]=16'h2ec5;
aud[6574]=16'h2eb6;
aud[6575]=16'h2ea7;
aud[6576]=16'h2e99;
aud[6577]=16'h2e8a;
aud[6578]=16'h2e7b;
aud[6579]=16'h2e6d;
aud[6580]=16'h2e5e;
aud[6581]=16'h2e4f;
aud[6582]=16'h2e40;
aud[6583]=16'h2e31;
aud[6584]=16'h2e22;
aud[6585]=16'h2e14;
aud[6586]=16'h2e05;
aud[6587]=16'h2df6;
aud[6588]=16'h2de7;
aud[6589]=16'h2dd8;
aud[6590]=16'h2dc9;
aud[6591]=16'h2dba;
aud[6592]=16'h2dab;
aud[6593]=16'h2d9c;
aud[6594]=16'h2d8d;
aud[6595]=16'h2d7e;
aud[6596]=16'h2d6f;
aud[6597]=16'h2d60;
aud[6598]=16'h2d50;
aud[6599]=16'h2d41;
aud[6600]=16'h2d32;
aud[6601]=16'h2d23;
aud[6602]=16'h2d14;
aud[6603]=16'h2d04;
aud[6604]=16'h2cf5;
aud[6605]=16'h2ce6;
aud[6606]=16'h2cd7;
aud[6607]=16'h2cc7;
aud[6608]=16'h2cb8;
aud[6609]=16'h2ca9;
aud[6610]=16'h2c99;
aud[6611]=16'h2c8a;
aud[6612]=16'h2c7a;
aud[6613]=16'h2c6b;
aud[6614]=16'h2c5c;
aud[6615]=16'h2c4c;
aud[6616]=16'h2c3d;
aud[6617]=16'h2c2d;
aud[6618]=16'h2c1e;
aud[6619]=16'h2c0e;
aud[6620]=16'h2bfe;
aud[6621]=16'h2bef;
aud[6622]=16'h2bdf;
aud[6623]=16'h2bd0;
aud[6624]=16'h2bc0;
aud[6625]=16'h2bb0;
aud[6626]=16'h2ba1;
aud[6627]=16'h2b91;
aud[6628]=16'h2b81;
aud[6629]=16'h2b71;
aud[6630]=16'h2b62;
aud[6631]=16'h2b52;
aud[6632]=16'h2b42;
aud[6633]=16'h2b32;
aud[6634]=16'h2b22;
aud[6635]=16'h2b13;
aud[6636]=16'h2b03;
aud[6637]=16'h2af3;
aud[6638]=16'h2ae3;
aud[6639]=16'h2ad3;
aud[6640]=16'h2ac3;
aud[6641]=16'h2ab3;
aud[6642]=16'h2aa3;
aud[6643]=16'h2a93;
aud[6644]=16'h2a83;
aud[6645]=16'h2a73;
aud[6646]=16'h2a63;
aud[6647]=16'h2a53;
aud[6648]=16'h2a43;
aud[6649]=16'h2a33;
aud[6650]=16'h2a23;
aud[6651]=16'h2a12;
aud[6652]=16'h2a02;
aud[6653]=16'h29f2;
aud[6654]=16'h29e2;
aud[6655]=16'h29d2;
aud[6656]=16'h29c1;
aud[6657]=16'h29b1;
aud[6658]=16'h29a1;
aud[6659]=16'h2991;
aud[6660]=16'h2980;
aud[6661]=16'h2970;
aud[6662]=16'h2960;
aud[6663]=16'h294f;
aud[6664]=16'h293f;
aud[6665]=16'h292e;
aud[6666]=16'h291e;
aud[6667]=16'h290e;
aud[6668]=16'h28fd;
aud[6669]=16'h28ed;
aud[6670]=16'h28dc;
aud[6671]=16'h28cc;
aud[6672]=16'h28bb;
aud[6673]=16'h28aa;
aud[6674]=16'h289a;
aud[6675]=16'h2889;
aud[6676]=16'h2879;
aud[6677]=16'h2868;
aud[6678]=16'h2857;
aud[6679]=16'h2847;
aud[6680]=16'h2836;
aud[6681]=16'h2825;
aud[6682]=16'h2815;
aud[6683]=16'h2804;
aud[6684]=16'h27f3;
aud[6685]=16'h27e2;
aud[6686]=16'h27d2;
aud[6687]=16'h27c1;
aud[6688]=16'h27b0;
aud[6689]=16'h279f;
aud[6690]=16'h278e;
aud[6691]=16'h277e;
aud[6692]=16'h276d;
aud[6693]=16'h275c;
aud[6694]=16'h274b;
aud[6695]=16'h273a;
aud[6696]=16'h2729;
aud[6697]=16'h2718;
aud[6698]=16'h2707;
aud[6699]=16'h26f6;
aud[6700]=16'h26e5;
aud[6701]=16'h26d4;
aud[6702]=16'h26c3;
aud[6703]=16'h26b2;
aud[6704]=16'h26a1;
aud[6705]=16'h2690;
aud[6706]=16'h267e;
aud[6707]=16'h266d;
aud[6708]=16'h265c;
aud[6709]=16'h264b;
aud[6710]=16'h263a;
aud[6711]=16'h2629;
aud[6712]=16'h2617;
aud[6713]=16'h2606;
aud[6714]=16'h25f5;
aud[6715]=16'h25e4;
aud[6716]=16'h25d2;
aud[6717]=16'h25c1;
aud[6718]=16'h25b0;
aud[6719]=16'h259e;
aud[6720]=16'h258d;
aud[6721]=16'h257c;
aud[6722]=16'h256a;
aud[6723]=16'h2559;
aud[6724]=16'h2547;
aud[6725]=16'h2536;
aud[6726]=16'h2524;
aud[6727]=16'h2513;
aud[6728]=16'h2501;
aud[6729]=16'h24f0;
aud[6730]=16'h24de;
aud[6731]=16'h24cd;
aud[6732]=16'h24bb;
aud[6733]=16'h24aa;
aud[6734]=16'h2498;
aud[6735]=16'h2487;
aud[6736]=16'h2475;
aud[6737]=16'h2463;
aud[6738]=16'h2452;
aud[6739]=16'h2440;
aud[6740]=16'h242e;
aud[6741]=16'h241d;
aud[6742]=16'h240b;
aud[6743]=16'h23f9;
aud[6744]=16'h23e7;
aud[6745]=16'h23d6;
aud[6746]=16'h23c4;
aud[6747]=16'h23b2;
aud[6748]=16'h23a0;
aud[6749]=16'h238e;
aud[6750]=16'h237d;
aud[6751]=16'h236b;
aud[6752]=16'h2359;
aud[6753]=16'h2347;
aud[6754]=16'h2335;
aud[6755]=16'h2323;
aud[6756]=16'h2311;
aud[6757]=16'h22ff;
aud[6758]=16'h22ed;
aud[6759]=16'h22db;
aud[6760]=16'h22c9;
aud[6761]=16'h22b7;
aud[6762]=16'h22a5;
aud[6763]=16'h2293;
aud[6764]=16'h2281;
aud[6765]=16'h226f;
aud[6766]=16'h225d;
aud[6767]=16'h224b;
aud[6768]=16'h2239;
aud[6769]=16'h2227;
aud[6770]=16'h2215;
aud[6771]=16'h2202;
aud[6772]=16'h21f0;
aud[6773]=16'h21de;
aud[6774]=16'h21cc;
aud[6775]=16'h21ba;
aud[6776]=16'h21a7;
aud[6777]=16'h2195;
aud[6778]=16'h2183;
aud[6779]=16'h2171;
aud[6780]=16'h215e;
aud[6781]=16'h214c;
aud[6782]=16'h213a;
aud[6783]=16'h2127;
aud[6784]=16'h2115;
aud[6785]=16'h2103;
aud[6786]=16'h20f0;
aud[6787]=16'h20de;
aud[6788]=16'h20cb;
aud[6789]=16'h20b9;
aud[6790]=16'h20a7;
aud[6791]=16'h2094;
aud[6792]=16'h2082;
aud[6793]=16'h206f;
aud[6794]=16'h205d;
aud[6795]=16'h204a;
aud[6796]=16'h2038;
aud[6797]=16'h2025;
aud[6798]=16'h2013;
aud[6799]=16'h2000;
aud[6800]=16'h1fed;
aud[6801]=16'h1fdb;
aud[6802]=16'h1fc8;
aud[6803]=16'h1fb6;
aud[6804]=16'h1fa3;
aud[6805]=16'h1f90;
aud[6806]=16'h1f7e;
aud[6807]=16'h1f6b;
aud[6808]=16'h1f58;
aud[6809]=16'h1f46;
aud[6810]=16'h1f33;
aud[6811]=16'h1f20;
aud[6812]=16'h1f0d;
aud[6813]=16'h1efb;
aud[6814]=16'h1ee8;
aud[6815]=16'h1ed5;
aud[6816]=16'h1ec2;
aud[6817]=16'h1eaf;
aud[6818]=16'h1e9d;
aud[6819]=16'h1e8a;
aud[6820]=16'h1e77;
aud[6821]=16'h1e64;
aud[6822]=16'h1e51;
aud[6823]=16'h1e3e;
aud[6824]=16'h1e2b;
aud[6825]=16'h1e18;
aud[6826]=16'h1e06;
aud[6827]=16'h1df3;
aud[6828]=16'h1de0;
aud[6829]=16'h1dcd;
aud[6830]=16'h1dba;
aud[6831]=16'h1da7;
aud[6832]=16'h1d94;
aud[6833]=16'h1d81;
aud[6834]=16'h1d6e;
aud[6835]=16'h1d5b;
aud[6836]=16'h1d47;
aud[6837]=16'h1d34;
aud[6838]=16'h1d21;
aud[6839]=16'h1d0e;
aud[6840]=16'h1cfb;
aud[6841]=16'h1ce8;
aud[6842]=16'h1cd5;
aud[6843]=16'h1cc2;
aud[6844]=16'h1cae;
aud[6845]=16'h1c9b;
aud[6846]=16'h1c88;
aud[6847]=16'h1c75;
aud[6848]=16'h1c62;
aud[6849]=16'h1c4e;
aud[6850]=16'h1c3b;
aud[6851]=16'h1c28;
aud[6852]=16'h1c15;
aud[6853]=16'h1c01;
aud[6854]=16'h1bee;
aud[6855]=16'h1bdb;
aud[6856]=16'h1bc8;
aud[6857]=16'h1bb4;
aud[6858]=16'h1ba1;
aud[6859]=16'h1b8d;
aud[6860]=16'h1b7a;
aud[6861]=16'h1b67;
aud[6862]=16'h1b53;
aud[6863]=16'h1b40;
aud[6864]=16'h1b2d;
aud[6865]=16'h1b19;
aud[6866]=16'h1b06;
aud[6867]=16'h1af2;
aud[6868]=16'h1adf;
aud[6869]=16'h1acb;
aud[6870]=16'h1ab8;
aud[6871]=16'h1aa4;
aud[6872]=16'h1a91;
aud[6873]=16'h1a7d;
aud[6874]=16'h1a6a;
aud[6875]=16'h1a56;
aud[6876]=16'h1a43;
aud[6877]=16'h1a2f;
aud[6878]=16'h1a1c;
aud[6879]=16'h1a08;
aud[6880]=16'h19f4;
aud[6881]=16'h19e1;
aud[6882]=16'h19cd;
aud[6883]=16'h19ba;
aud[6884]=16'h19a6;
aud[6885]=16'h1992;
aud[6886]=16'h197f;
aud[6887]=16'h196b;
aud[6888]=16'h1957;
aud[6889]=16'h1943;
aud[6890]=16'h1930;
aud[6891]=16'h191c;
aud[6892]=16'h1908;
aud[6893]=16'h18f5;
aud[6894]=16'h18e1;
aud[6895]=16'h18cd;
aud[6896]=16'h18b9;
aud[6897]=16'h18a5;
aud[6898]=16'h1892;
aud[6899]=16'h187e;
aud[6900]=16'h186a;
aud[6901]=16'h1856;
aud[6902]=16'h1842;
aud[6903]=16'h182f;
aud[6904]=16'h181b;
aud[6905]=16'h1807;
aud[6906]=16'h17f3;
aud[6907]=16'h17df;
aud[6908]=16'h17cb;
aud[6909]=16'h17b7;
aud[6910]=16'h17a3;
aud[6911]=16'h178f;
aud[6912]=16'h177b;
aud[6913]=16'h1767;
aud[6914]=16'h1753;
aud[6915]=16'h1740;
aud[6916]=16'h172c;
aud[6917]=16'h1718;
aud[6918]=16'h1704;
aud[6919]=16'h16f0;
aud[6920]=16'h16db;
aud[6921]=16'h16c7;
aud[6922]=16'h16b3;
aud[6923]=16'h169f;
aud[6924]=16'h168b;
aud[6925]=16'h1677;
aud[6926]=16'h1663;
aud[6927]=16'h164f;
aud[6928]=16'h163b;
aud[6929]=16'h1627;
aud[6930]=16'h1613;
aud[6931]=16'h15ff;
aud[6932]=16'h15ea;
aud[6933]=16'h15d6;
aud[6934]=16'h15c2;
aud[6935]=16'h15ae;
aud[6936]=16'h159a;
aud[6937]=16'h1586;
aud[6938]=16'h1571;
aud[6939]=16'h155d;
aud[6940]=16'h1549;
aud[6941]=16'h1535;
aud[6942]=16'h1520;
aud[6943]=16'h150c;
aud[6944]=16'h14f8;
aud[6945]=16'h14e4;
aud[6946]=16'h14cf;
aud[6947]=16'h14bb;
aud[6948]=16'h14a7;
aud[6949]=16'h1492;
aud[6950]=16'h147e;
aud[6951]=16'h146a;
aud[6952]=16'h1455;
aud[6953]=16'h1441;
aud[6954]=16'h142d;
aud[6955]=16'h1418;
aud[6956]=16'h1404;
aud[6957]=16'h13f0;
aud[6958]=16'h13db;
aud[6959]=16'h13c7;
aud[6960]=16'h13b3;
aud[6961]=16'h139e;
aud[6962]=16'h138a;
aud[6963]=16'h1375;
aud[6964]=16'h1361;
aud[6965]=16'h134c;
aud[6966]=16'h1338;
aud[6967]=16'h1323;
aud[6968]=16'h130f;
aud[6969]=16'h12fb;
aud[6970]=16'h12e6;
aud[6971]=16'h12d2;
aud[6972]=16'h12bd;
aud[6973]=16'h12a9;
aud[6974]=16'h1294;
aud[6975]=16'h127f;
aud[6976]=16'h126b;
aud[6977]=16'h1256;
aud[6978]=16'h1242;
aud[6979]=16'h122d;
aud[6980]=16'h1219;
aud[6981]=16'h1204;
aud[6982]=16'h11f0;
aud[6983]=16'h11db;
aud[6984]=16'h11c6;
aud[6985]=16'h11b2;
aud[6986]=16'h119d;
aud[6987]=16'h1189;
aud[6988]=16'h1174;
aud[6989]=16'h115f;
aud[6990]=16'h114b;
aud[6991]=16'h1136;
aud[6992]=16'h1121;
aud[6993]=16'h110d;
aud[6994]=16'h10f8;
aud[6995]=16'h10e3;
aud[6996]=16'h10cf;
aud[6997]=16'h10ba;
aud[6998]=16'h10a5;
aud[6999]=16'h1090;
aud[7000]=16'h107c;
aud[7001]=16'h1067;
aud[7002]=16'h1052;
aud[7003]=16'h103e;
aud[7004]=16'h1029;
aud[7005]=16'h1014;
aud[7006]=16'hfff;
aud[7007]=16'hfeb;
aud[7008]=16'hfd6;
aud[7009]=16'hfc1;
aud[7010]=16'hfac;
aud[7011]=16'hf97;
aud[7012]=16'hf83;
aud[7013]=16'hf6e;
aud[7014]=16'hf59;
aud[7015]=16'hf44;
aud[7016]=16'hf2f;
aud[7017]=16'hf1a;
aud[7018]=16'hf06;
aud[7019]=16'hef1;
aud[7020]=16'hedc;
aud[7021]=16'hec7;
aud[7022]=16'heb2;
aud[7023]=16'he9d;
aud[7024]=16'he88;
aud[7025]=16'he74;
aud[7026]=16'he5f;
aud[7027]=16'he4a;
aud[7028]=16'he35;
aud[7029]=16'he20;
aud[7030]=16'he0b;
aud[7031]=16'hdf6;
aud[7032]=16'hde1;
aud[7033]=16'hdcc;
aud[7034]=16'hdb7;
aud[7035]=16'hda2;
aud[7036]=16'hd8d;
aud[7037]=16'hd78;
aud[7038]=16'hd63;
aud[7039]=16'hd4e;
aud[7040]=16'hd39;
aud[7041]=16'hd24;
aud[7042]=16'hd0f;
aud[7043]=16'hcfa;
aud[7044]=16'hce5;
aud[7045]=16'hcd0;
aud[7046]=16'hcbb;
aud[7047]=16'hca6;
aud[7048]=16'hc91;
aud[7049]=16'hc7c;
aud[7050]=16'hc67;
aud[7051]=16'hc52;
aud[7052]=16'hc3d;
aud[7053]=16'hc28;
aud[7054]=16'hc13;
aud[7055]=16'hbfe;
aud[7056]=16'hbe9;
aud[7057]=16'hbd4;
aud[7058]=16'hbbf;
aud[7059]=16'hbaa;
aud[7060]=16'hb95;
aud[7061]=16'hb80;
aud[7062]=16'hb6a;
aud[7063]=16'hb55;
aud[7064]=16'hb40;
aud[7065]=16'hb2b;
aud[7066]=16'hb16;
aud[7067]=16'hb01;
aud[7068]=16'haec;
aud[7069]=16'had7;
aud[7070]=16'hac1;
aud[7071]=16'haac;
aud[7072]=16'ha97;
aud[7073]=16'ha82;
aud[7074]=16'ha6d;
aud[7075]=16'ha58;
aud[7076]=16'ha43;
aud[7077]=16'ha2d;
aud[7078]=16'ha18;
aud[7079]=16'ha03;
aud[7080]=16'h9ee;
aud[7081]=16'h9d9;
aud[7082]=16'h9c3;
aud[7083]=16'h9ae;
aud[7084]=16'h999;
aud[7085]=16'h984;
aud[7086]=16'h96f;
aud[7087]=16'h959;
aud[7088]=16'h944;
aud[7089]=16'h92f;
aud[7090]=16'h91a;
aud[7091]=16'h905;
aud[7092]=16'h8ef;
aud[7093]=16'h8da;
aud[7094]=16'h8c5;
aud[7095]=16'h8b0;
aud[7096]=16'h89a;
aud[7097]=16'h885;
aud[7098]=16'h870;
aud[7099]=16'h85b;
aud[7100]=16'h845;
aud[7101]=16'h830;
aud[7102]=16'h81b;
aud[7103]=16'h805;
aud[7104]=16'h7f0;
aud[7105]=16'h7db;
aud[7106]=16'h7c6;
aud[7107]=16'h7b0;
aud[7108]=16'h79b;
aud[7109]=16'h786;
aud[7110]=16'h770;
aud[7111]=16'h75b;
aud[7112]=16'h746;
aud[7113]=16'h731;
aud[7114]=16'h71b;
aud[7115]=16'h706;
aud[7116]=16'h6f1;
aud[7117]=16'h6db;
aud[7118]=16'h6c6;
aud[7119]=16'h6b1;
aud[7120]=16'h69b;
aud[7121]=16'h686;
aud[7122]=16'h671;
aud[7123]=16'h65b;
aud[7124]=16'h646;
aud[7125]=16'h631;
aud[7126]=16'h61b;
aud[7127]=16'h606;
aud[7128]=16'h5f1;
aud[7129]=16'h5db;
aud[7130]=16'h5c6;
aud[7131]=16'h5b0;
aud[7132]=16'h59b;
aud[7133]=16'h586;
aud[7134]=16'h570;
aud[7135]=16'h55b;
aud[7136]=16'h546;
aud[7137]=16'h530;
aud[7138]=16'h51b;
aud[7139]=16'h505;
aud[7140]=16'h4f0;
aud[7141]=16'h4db;
aud[7142]=16'h4c5;
aud[7143]=16'h4b0;
aud[7144]=16'h49b;
aud[7145]=16'h485;
aud[7146]=16'h470;
aud[7147]=16'h45a;
aud[7148]=16'h445;
aud[7149]=16'h430;
aud[7150]=16'h41a;
aud[7151]=16'h405;
aud[7152]=16'h3ef;
aud[7153]=16'h3da;
aud[7154]=16'h3c5;
aud[7155]=16'h3af;
aud[7156]=16'h39a;
aud[7157]=16'h384;
aud[7158]=16'h36f;
aud[7159]=16'h359;
aud[7160]=16'h344;
aud[7161]=16'h32f;
aud[7162]=16'h319;
aud[7163]=16'h304;
aud[7164]=16'h2ee;
aud[7165]=16'h2d9;
aud[7166]=16'h2c4;
aud[7167]=16'h2ae;
aud[7168]=16'h299;
aud[7169]=16'h283;
aud[7170]=16'h26e;
aud[7171]=16'h258;
aud[7172]=16'h243;
aud[7173]=16'h22e;
aud[7174]=16'h218;
aud[7175]=16'h203;
aud[7176]=16'h1ed;
aud[7177]=16'h1d8;
aud[7178]=16'h1c2;
aud[7179]=16'h1ad;
aud[7180]=16'h197;
aud[7181]=16'h182;
aud[7182]=16'h16d;
aud[7183]=16'h157;
aud[7184]=16'h142;
aud[7185]=16'h12c;
aud[7186]=16'h117;
aud[7187]=16'h101;
aud[7188]=16'hec;
aud[7189]=16'hd6;
aud[7190]=16'hc1;
aud[7191]=16'hac;
aud[7192]=16'h96;
aud[7193]=16'h81;
aud[7194]=16'h6b;
aud[7195]=16'h56;
aud[7196]=16'h40;
aud[7197]=16'h2b;
aud[7198]=16'h15;
aud[7199]=16'h0;
aud[7200]=16'hffeb;
aud[7201]=16'hffd5;
aud[7202]=16'hffc0;
aud[7203]=16'hffaa;
aud[7204]=16'hff95;
aud[7205]=16'hff7f;
aud[7206]=16'hff6a;
aud[7207]=16'hff54;
aud[7208]=16'hff3f;
aud[7209]=16'hff2a;
aud[7210]=16'hff14;
aud[7211]=16'hfeff;
aud[7212]=16'hfee9;
aud[7213]=16'hfed4;
aud[7214]=16'hfebe;
aud[7215]=16'hfea9;
aud[7216]=16'hfe93;
aud[7217]=16'hfe7e;
aud[7218]=16'hfe69;
aud[7219]=16'hfe53;
aud[7220]=16'hfe3e;
aud[7221]=16'hfe28;
aud[7222]=16'hfe13;
aud[7223]=16'hfdfd;
aud[7224]=16'hfde8;
aud[7225]=16'hfdd2;
aud[7226]=16'hfdbd;
aud[7227]=16'hfda8;
aud[7228]=16'hfd92;
aud[7229]=16'hfd7d;
aud[7230]=16'hfd67;
aud[7231]=16'hfd52;
aud[7232]=16'hfd3c;
aud[7233]=16'hfd27;
aud[7234]=16'hfd12;
aud[7235]=16'hfcfc;
aud[7236]=16'hfce7;
aud[7237]=16'hfcd1;
aud[7238]=16'hfcbc;
aud[7239]=16'hfca7;
aud[7240]=16'hfc91;
aud[7241]=16'hfc7c;
aud[7242]=16'hfc66;
aud[7243]=16'hfc51;
aud[7244]=16'hfc3b;
aud[7245]=16'hfc26;
aud[7246]=16'hfc11;
aud[7247]=16'hfbfb;
aud[7248]=16'hfbe6;
aud[7249]=16'hfbd0;
aud[7250]=16'hfbbb;
aud[7251]=16'hfba6;
aud[7252]=16'hfb90;
aud[7253]=16'hfb7b;
aud[7254]=16'hfb65;
aud[7255]=16'hfb50;
aud[7256]=16'hfb3b;
aud[7257]=16'hfb25;
aud[7258]=16'hfb10;
aud[7259]=16'hfafb;
aud[7260]=16'hfae5;
aud[7261]=16'hfad0;
aud[7262]=16'hfaba;
aud[7263]=16'hfaa5;
aud[7264]=16'hfa90;
aud[7265]=16'hfa7a;
aud[7266]=16'hfa65;
aud[7267]=16'hfa50;
aud[7268]=16'hfa3a;
aud[7269]=16'hfa25;
aud[7270]=16'hfa0f;
aud[7271]=16'hf9fa;
aud[7272]=16'hf9e5;
aud[7273]=16'hf9cf;
aud[7274]=16'hf9ba;
aud[7275]=16'hf9a5;
aud[7276]=16'hf98f;
aud[7277]=16'hf97a;
aud[7278]=16'hf965;
aud[7279]=16'hf94f;
aud[7280]=16'hf93a;
aud[7281]=16'hf925;
aud[7282]=16'hf90f;
aud[7283]=16'hf8fa;
aud[7284]=16'hf8e5;
aud[7285]=16'hf8cf;
aud[7286]=16'hf8ba;
aud[7287]=16'hf8a5;
aud[7288]=16'hf890;
aud[7289]=16'hf87a;
aud[7290]=16'hf865;
aud[7291]=16'hf850;
aud[7292]=16'hf83a;
aud[7293]=16'hf825;
aud[7294]=16'hf810;
aud[7295]=16'hf7fb;
aud[7296]=16'hf7e5;
aud[7297]=16'hf7d0;
aud[7298]=16'hf7bb;
aud[7299]=16'hf7a5;
aud[7300]=16'hf790;
aud[7301]=16'hf77b;
aud[7302]=16'hf766;
aud[7303]=16'hf750;
aud[7304]=16'hf73b;
aud[7305]=16'hf726;
aud[7306]=16'hf711;
aud[7307]=16'hf6fb;
aud[7308]=16'hf6e6;
aud[7309]=16'hf6d1;
aud[7310]=16'hf6bc;
aud[7311]=16'hf6a7;
aud[7312]=16'hf691;
aud[7313]=16'hf67c;
aud[7314]=16'hf667;
aud[7315]=16'hf652;
aud[7316]=16'hf63d;
aud[7317]=16'hf627;
aud[7318]=16'hf612;
aud[7319]=16'hf5fd;
aud[7320]=16'hf5e8;
aud[7321]=16'hf5d3;
aud[7322]=16'hf5bd;
aud[7323]=16'hf5a8;
aud[7324]=16'hf593;
aud[7325]=16'hf57e;
aud[7326]=16'hf569;
aud[7327]=16'hf554;
aud[7328]=16'hf53f;
aud[7329]=16'hf529;
aud[7330]=16'hf514;
aud[7331]=16'hf4ff;
aud[7332]=16'hf4ea;
aud[7333]=16'hf4d5;
aud[7334]=16'hf4c0;
aud[7335]=16'hf4ab;
aud[7336]=16'hf496;
aud[7337]=16'hf480;
aud[7338]=16'hf46b;
aud[7339]=16'hf456;
aud[7340]=16'hf441;
aud[7341]=16'hf42c;
aud[7342]=16'hf417;
aud[7343]=16'hf402;
aud[7344]=16'hf3ed;
aud[7345]=16'hf3d8;
aud[7346]=16'hf3c3;
aud[7347]=16'hf3ae;
aud[7348]=16'hf399;
aud[7349]=16'hf384;
aud[7350]=16'hf36f;
aud[7351]=16'hf35a;
aud[7352]=16'hf345;
aud[7353]=16'hf330;
aud[7354]=16'hf31b;
aud[7355]=16'hf306;
aud[7356]=16'hf2f1;
aud[7357]=16'hf2dc;
aud[7358]=16'hf2c7;
aud[7359]=16'hf2b2;
aud[7360]=16'hf29d;
aud[7361]=16'hf288;
aud[7362]=16'hf273;
aud[7363]=16'hf25e;
aud[7364]=16'hf249;
aud[7365]=16'hf234;
aud[7366]=16'hf21f;
aud[7367]=16'hf20a;
aud[7368]=16'hf1f5;
aud[7369]=16'hf1e0;
aud[7370]=16'hf1cb;
aud[7371]=16'hf1b6;
aud[7372]=16'hf1a1;
aud[7373]=16'hf18c;
aud[7374]=16'hf178;
aud[7375]=16'hf163;
aud[7376]=16'hf14e;
aud[7377]=16'hf139;
aud[7378]=16'hf124;
aud[7379]=16'hf10f;
aud[7380]=16'hf0fa;
aud[7381]=16'hf0e6;
aud[7382]=16'hf0d1;
aud[7383]=16'hf0bc;
aud[7384]=16'hf0a7;
aud[7385]=16'hf092;
aud[7386]=16'hf07d;
aud[7387]=16'hf069;
aud[7388]=16'hf054;
aud[7389]=16'hf03f;
aud[7390]=16'hf02a;
aud[7391]=16'hf015;
aud[7392]=16'hf001;
aud[7393]=16'hefec;
aud[7394]=16'hefd7;
aud[7395]=16'hefc2;
aud[7396]=16'hefae;
aud[7397]=16'hef99;
aud[7398]=16'hef84;
aud[7399]=16'hef70;
aud[7400]=16'hef5b;
aud[7401]=16'hef46;
aud[7402]=16'hef31;
aud[7403]=16'hef1d;
aud[7404]=16'hef08;
aud[7405]=16'heef3;
aud[7406]=16'heedf;
aud[7407]=16'heeca;
aud[7408]=16'heeb5;
aud[7409]=16'heea1;
aud[7410]=16'hee8c;
aud[7411]=16'hee77;
aud[7412]=16'hee63;
aud[7413]=16'hee4e;
aud[7414]=16'hee3a;
aud[7415]=16'hee25;
aud[7416]=16'hee10;
aud[7417]=16'hedfc;
aud[7418]=16'hede7;
aud[7419]=16'hedd3;
aud[7420]=16'hedbe;
aud[7421]=16'hedaa;
aud[7422]=16'hed95;
aud[7423]=16'hed81;
aud[7424]=16'hed6c;
aud[7425]=16'hed57;
aud[7426]=16'hed43;
aud[7427]=16'hed2e;
aud[7428]=16'hed1a;
aud[7429]=16'hed05;
aud[7430]=16'hecf1;
aud[7431]=16'hecdd;
aud[7432]=16'hecc8;
aud[7433]=16'hecb4;
aud[7434]=16'hec9f;
aud[7435]=16'hec8b;
aud[7436]=16'hec76;
aud[7437]=16'hec62;
aud[7438]=16'hec4d;
aud[7439]=16'hec39;
aud[7440]=16'hec25;
aud[7441]=16'hec10;
aud[7442]=16'hebfc;
aud[7443]=16'hebe8;
aud[7444]=16'hebd3;
aud[7445]=16'hebbf;
aud[7446]=16'hebab;
aud[7447]=16'heb96;
aud[7448]=16'heb82;
aud[7449]=16'heb6e;
aud[7450]=16'heb59;
aud[7451]=16'heb45;
aud[7452]=16'heb31;
aud[7453]=16'heb1c;
aud[7454]=16'heb08;
aud[7455]=16'heaf4;
aud[7456]=16'heae0;
aud[7457]=16'heacb;
aud[7458]=16'heab7;
aud[7459]=16'heaa3;
aud[7460]=16'hea8f;
aud[7461]=16'hea7a;
aud[7462]=16'hea66;
aud[7463]=16'hea52;
aud[7464]=16'hea3e;
aud[7465]=16'hea2a;
aud[7466]=16'hea16;
aud[7467]=16'hea01;
aud[7468]=16'he9ed;
aud[7469]=16'he9d9;
aud[7470]=16'he9c5;
aud[7471]=16'he9b1;
aud[7472]=16'he99d;
aud[7473]=16'he989;
aud[7474]=16'he975;
aud[7475]=16'he961;
aud[7476]=16'he94d;
aud[7477]=16'he939;
aud[7478]=16'he925;
aud[7479]=16'he910;
aud[7480]=16'he8fc;
aud[7481]=16'he8e8;
aud[7482]=16'he8d4;
aud[7483]=16'he8c0;
aud[7484]=16'he8ad;
aud[7485]=16'he899;
aud[7486]=16'he885;
aud[7487]=16'he871;
aud[7488]=16'he85d;
aud[7489]=16'he849;
aud[7490]=16'he835;
aud[7491]=16'he821;
aud[7492]=16'he80d;
aud[7493]=16'he7f9;
aud[7494]=16'he7e5;
aud[7495]=16'he7d1;
aud[7496]=16'he7be;
aud[7497]=16'he7aa;
aud[7498]=16'he796;
aud[7499]=16'he782;
aud[7500]=16'he76e;
aud[7501]=16'he75b;
aud[7502]=16'he747;
aud[7503]=16'he733;
aud[7504]=16'he71f;
aud[7505]=16'he70b;
aud[7506]=16'he6f8;
aud[7507]=16'he6e4;
aud[7508]=16'he6d0;
aud[7509]=16'he6bd;
aud[7510]=16'he6a9;
aud[7511]=16'he695;
aud[7512]=16'he681;
aud[7513]=16'he66e;
aud[7514]=16'he65a;
aud[7515]=16'he646;
aud[7516]=16'he633;
aud[7517]=16'he61f;
aud[7518]=16'he60c;
aud[7519]=16'he5f8;
aud[7520]=16'he5e4;
aud[7521]=16'he5d1;
aud[7522]=16'he5bd;
aud[7523]=16'he5aa;
aud[7524]=16'he596;
aud[7525]=16'he583;
aud[7526]=16'he56f;
aud[7527]=16'he55c;
aud[7528]=16'he548;
aud[7529]=16'he535;
aud[7530]=16'he521;
aud[7531]=16'he50e;
aud[7532]=16'he4fa;
aud[7533]=16'he4e7;
aud[7534]=16'he4d3;
aud[7535]=16'he4c0;
aud[7536]=16'he4ad;
aud[7537]=16'he499;
aud[7538]=16'he486;
aud[7539]=16'he473;
aud[7540]=16'he45f;
aud[7541]=16'he44c;
aud[7542]=16'he438;
aud[7543]=16'he425;
aud[7544]=16'he412;
aud[7545]=16'he3ff;
aud[7546]=16'he3eb;
aud[7547]=16'he3d8;
aud[7548]=16'he3c5;
aud[7549]=16'he3b2;
aud[7550]=16'he39e;
aud[7551]=16'he38b;
aud[7552]=16'he378;
aud[7553]=16'he365;
aud[7554]=16'he352;
aud[7555]=16'he33e;
aud[7556]=16'he32b;
aud[7557]=16'he318;
aud[7558]=16'he305;
aud[7559]=16'he2f2;
aud[7560]=16'he2df;
aud[7561]=16'he2cc;
aud[7562]=16'he2b9;
aud[7563]=16'he2a5;
aud[7564]=16'he292;
aud[7565]=16'he27f;
aud[7566]=16'he26c;
aud[7567]=16'he259;
aud[7568]=16'he246;
aud[7569]=16'he233;
aud[7570]=16'he220;
aud[7571]=16'he20d;
aud[7572]=16'he1fa;
aud[7573]=16'he1e8;
aud[7574]=16'he1d5;
aud[7575]=16'he1c2;
aud[7576]=16'he1af;
aud[7577]=16'he19c;
aud[7578]=16'he189;
aud[7579]=16'he176;
aud[7580]=16'he163;
aud[7581]=16'he151;
aud[7582]=16'he13e;
aud[7583]=16'he12b;
aud[7584]=16'he118;
aud[7585]=16'he105;
aud[7586]=16'he0f3;
aud[7587]=16'he0e0;
aud[7588]=16'he0cd;
aud[7589]=16'he0ba;
aud[7590]=16'he0a8;
aud[7591]=16'he095;
aud[7592]=16'he082;
aud[7593]=16'he070;
aud[7594]=16'he05d;
aud[7595]=16'he04a;
aud[7596]=16'he038;
aud[7597]=16'he025;
aud[7598]=16'he013;
aud[7599]=16'he000;
aud[7600]=16'hdfed;
aud[7601]=16'hdfdb;
aud[7602]=16'hdfc8;
aud[7603]=16'hdfb6;
aud[7604]=16'hdfa3;
aud[7605]=16'hdf91;
aud[7606]=16'hdf7e;
aud[7607]=16'hdf6c;
aud[7608]=16'hdf59;
aud[7609]=16'hdf47;
aud[7610]=16'hdf35;
aud[7611]=16'hdf22;
aud[7612]=16'hdf10;
aud[7613]=16'hdefd;
aud[7614]=16'hdeeb;
aud[7615]=16'hded9;
aud[7616]=16'hdec6;
aud[7617]=16'hdeb4;
aud[7618]=16'hdea2;
aud[7619]=16'hde8f;
aud[7620]=16'hde7d;
aud[7621]=16'hde6b;
aud[7622]=16'hde59;
aud[7623]=16'hde46;
aud[7624]=16'hde34;
aud[7625]=16'hde22;
aud[7626]=16'hde10;
aud[7627]=16'hddfe;
aud[7628]=16'hddeb;
aud[7629]=16'hddd9;
aud[7630]=16'hddc7;
aud[7631]=16'hddb5;
aud[7632]=16'hdda3;
aud[7633]=16'hdd91;
aud[7634]=16'hdd7f;
aud[7635]=16'hdd6d;
aud[7636]=16'hdd5b;
aud[7637]=16'hdd49;
aud[7638]=16'hdd37;
aud[7639]=16'hdd25;
aud[7640]=16'hdd13;
aud[7641]=16'hdd01;
aud[7642]=16'hdcef;
aud[7643]=16'hdcdd;
aud[7644]=16'hdccb;
aud[7645]=16'hdcb9;
aud[7646]=16'hdca7;
aud[7647]=16'hdc95;
aud[7648]=16'hdc83;
aud[7649]=16'hdc72;
aud[7650]=16'hdc60;
aud[7651]=16'hdc4e;
aud[7652]=16'hdc3c;
aud[7653]=16'hdc2a;
aud[7654]=16'hdc19;
aud[7655]=16'hdc07;
aud[7656]=16'hdbf5;
aud[7657]=16'hdbe3;
aud[7658]=16'hdbd2;
aud[7659]=16'hdbc0;
aud[7660]=16'hdbae;
aud[7661]=16'hdb9d;
aud[7662]=16'hdb8b;
aud[7663]=16'hdb79;
aud[7664]=16'hdb68;
aud[7665]=16'hdb56;
aud[7666]=16'hdb45;
aud[7667]=16'hdb33;
aud[7668]=16'hdb22;
aud[7669]=16'hdb10;
aud[7670]=16'hdaff;
aud[7671]=16'hdaed;
aud[7672]=16'hdadc;
aud[7673]=16'hdaca;
aud[7674]=16'hdab9;
aud[7675]=16'hdaa7;
aud[7676]=16'hda96;
aud[7677]=16'hda84;
aud[7678]=16'hda73;
aud[7679]=16'hda62;
aud[7680]=16'hda50;
aud[7681]=16'hda3f;
aud[7682]=16'hda2e;
aud[7683]=16'hda1c;
aud[7684]=16'hda0b;
aud[7685]=16'hd9fa;
aud[7686]=16'hd9e9;
aud[7687]=16'hd9d7;
aud[7688]=16'hd9c6;
aud[7689]=16'hd9b5;
aud[7690]=16'hd9a4;
aud[7691]=16'hd993;
aud[7692]=16'hd982;
aud[7693]=16'hd970;
aud[7694]=16'hd95f;
aud[7695]=16'hd94e;
aud[7696]=16'hd93d;
aud[7697]=16'hd92c;
aud[7698]=16'hd91b;
aud[7699]=16'hd90a;
aud[7700]=16'hd8f9;
aud[7701]=16'hd8e8;
aud[7702]=16'hd8d7;
aud[7703]=16'hd8c6;
aud[7704]=16'hd8b5;
aud[7705]=16'hd8a4;
aud[7706]=16'hd893;
aud[7707]=16'hd882;
aud[7708]=16'hd872;
aud[7709]=16'hd861;
aud[7710]=16'hd850;
aud[7711]=16'hd83f;
aud[7712]=16'hd82e;
aud[7713]=16'hd81e;
aud[7714]=16'hd80d;
aud[7715]=16'hd7fc;
aud[7716]=16'hd7eb;
aud[7717]=16'hd7db;
aud[7718]=16'hd7ca;
aud[7719]=16'hd7b9;
aud[7720]=16'hd7a9;
aud[7721]=16'hd798;
aud[7722]=16'hd787;
aud[7723]=16'hd777;
aud[7724]=16'hd766;
aud[7725]=16'hd756;
aud[7726]=16'hd745;
aud[7727]=16'hd734;
aud[7728]=16'hd724;
aud[7729]=16'hd713;
aud[7730]=16'hd703;
aud[7731]=16'hd6f2;
aud[7732]=16'hd6e2;
aud[7733]=16'hd6d2;
aud[7734]=16'hd6c1;
aud[7735]=16'hd6b1;
aud[7736]=16'hd6a0;
aud[7737]=16'hd690;
aud[7738]=16'hd680;
aud[7739]=16'hd66f;
aud[7740]=16'hd65f;
aud[7741]=16'hd64f;
aud[7742]=16'hd63f;
aud[7743]=16'hd62e;
aud[7744]=16'hd61e;
aud[7745]=16'hd60e;
aud[7746]=16'hd5fe;
aud[7747]=16'hd5ee;
aud[7748]=16'hd5dd;
aud[7749]=16'hd5cd;
aud[7750]=16'hd5bd;
aud[7751]=16'hd5ad;
aud[7752]=16'hd59d;
aud[7753]=16'hd58d;
aud[7754]=16'hd57d;
aud[7755]=16'hd56d;
aud[7756]=16'hd55d;
aud[7757]=16'hd54d;
aud[7758]=16'hd53d;
aud[7759]=16'hd52d;
aud[7760]=16'hd51d;
aud[7761]=16'hd50d;
aud[7762]=16'hd4fd;
aud[7763]=16'hd4ed;
aud[7764]=16'hd4de;
aud[7765]=16'hd4ce;
aud[7766]=16'hd4be;
aud[7767]=16'hd4ae;
aud[7768]=16'hd49e;
aud[7769]=16'hd48f;
aud[7770]=16'hd47f;
aud[7771]=16'hd46f;
aud[7772]=16'hd45f;
aud[7773]=16'hd450;
aud[7774]=16'hd440;
aud[7775]=16'hd430;
aud[7776]=16'hd421;
aud[7777]=16'hd411;
aud[7778]=16'hd402;
aud[7779]=16'hd3f2;
aud[7780]=16'hd3e2;
aud[7781]=16'hd3d3;
aud[7782]=16'hd3c3;
aud[7783]=16'hd3b4;
aud[7784]=16'hd3a4;
aud[7785]=16'hd395;
aud[7786]=16'hd386;
aud[7787]=16'hd376;
aud[7788]=16'hd367;
aud[7789]=16'hd357;
aud[7790]=16'hd348;
aud[7791]=16'hd339;
aud[7792]=16'hd329;
aud[7793]=16'hd31a;
aud[7794]=16'hd30b;
aud[7795]=16'hd2fc;
aud[7796]=16'hd2ec;
aud[7797]=16'hd2dd;
aud[7798]=16'hd2ce;
aud[7799]=16'hd2bf;
aud[7800]=16'hd2b0;
aud[7801]=16'hd2a0;
aud[7802]=16'hd291;
aud[7803]=16'hd282;
aud[7804]=16'hd273;
aud[7805]=16'hd264;
aud[7806]=16'hd255;
aud[7807]=16'hd246;
aud[7808]=16'hd237;
aud[7809]=16'hd228;
aud[7810]=16'hd219;
aud[7811]=16'hd20a;
aud[7812]=16'hd1fb;
aud[7813]=16'hd1ec;
aud[7814]=16'hd1de;
aud[7815]=16'hd1cf;
aud[7816]=16'hd1c0;
aud[7817]=16'hd1b1;
aud[7818]=16'hd1a2;
aud[7819]=16'hd193;
aud[7820]=16'hd185;
aud[7821]=16'hd176;
aud[7822]=16'hd167;
aud[7823]=16'hd159;
aud[7824]=16'hd14a;
aud[7825]=16'hd13b;
aud[7826]=16'hd12d;
aud[7827]=16'hd11e;
aud[7828]=16'hd10f;
aud[7829]=16'hd101;
aud[7830]=16'hd0f2;
aud[7831]=16'hd0e4;
aud[7832]=16'hd0d5;
aud[7833]=16'hd0c7;
aud[7834]=16'hd0b8;
aud[7835]=16'hd0aa;
aud[7836]=16'hd09b;
aud[7837]=16'hd08d;
aud[7838]=16'hd07f;
aud[7839]=16'hd070;
aud[7840]=16'hd062;
aud[7841]=16'hd054;
aud[7842]=16'hd045;
aud[7843]=16'hd037;
aud[7844]=16'hd029;
aud[7845]=16'hd01b;
aud[7846]=16'hd00c;
aud[7847]=16'hcffe;
aud[7848]=16'hcff0;
aud[7849]=16'hcfe2;
aud[7850]=16'hcfd4;
aud[7851]=16'hcfc6;
aud[7852]=16'hcfb8;
aud[7853]=16'hcfa9;
aud[7854]=16'hcf9b;
aud[7855]=16'hcf8d;
aud[7856]=16'hcf7f;
aud[7857]=16'hcf71;
aud[7858]=16'hcf63;
aud[7859]=16'hcf56;
aud[7860]=16'hcf48;
aud[7861]=16'hcf3a;
aud[7862]=16'hcf2c;
aud[7863]=16'hcf1e;
aud[7864]=16'hcf10;
aud[7865]=16'hcf02;
aud[7866]=16'hcef5;
aud[7867]=16'hcee7;
aud[7868]=16'hced9;
aud[7869]=16'hcecb;
aud[7870]=16'hcebe;
aud[7871]=16'hceb0;
aud[7872]=16'hcea2;
aud[7873]=16'hce95;
aud[7874]=16'hce87;
aud[7875]=16'hce79;
aud[7876]=16'hce6c;
aud[7877]=16'hce5e;
aud[7878]=16'hce51;
aud[7879]=16'hce43;
aud[7880]=16'hce36;
aud[7881]=16'hce28;
aud[7882]=16'hce1b;
aud[7883]=16'hce0d;
aud[7884]=16'hce00;
aud[7885]=16'hcdf3;
aud[7886]=16'hcde5;
aud[7887]=16'hcdd8;
aud[7888]=16'hcdcb;
aud[7889]=16'hcdbd;
aud[7890]=16'hcdb0;
aud[7891]=16'hcda3;
aud[7892]=16'hcd96;
aud[7893]=16'hcd88;
aud[7894]=16'hcd7b;
aud[7895]=16'hcd6e;
aud[7896]=16'hcd61;
aud[7897]=16'hcd54;
aud[7898]=16'hcd47;
aud[7899]=16'hcd3a;
aud[7900]=16'hcd2d;
aud[7901]=16'hcd20;
aud[7902]=16'hcd13;
aud[7903]=16'hcd06;
aud[7904]=16'hccf9;
aud[7905]=16'hccec;
aud[7906]=16'hccdf;
aud[7907]=16'hccd2;
aud[7908]=16'hccc5;
aud[7909]=16'hccb8;
aud[7910]=16'hccab;
aud[7911]=16'hcc9f;
aud[7912]=16'hcc92;
aud[7913]=16'hcc85;
aud[7914]=16'hcc78;
aud[7915]=16'hcc6c;
aud[7916]=16'hcc5f;
aud[7917]=16'hcc52;
aud[7918]=16'hcc46;
aud[7919]=16'hcc39;
aud[7920]=16'hcc2c;
aud[7921]=16'hcc20;
aud[7922]=16'hcc13;
aud[7923]=16'hcc07;
aud[7924]=16'hcbfa;
aud[7925]=16'hcbee;
aud[7926]=16'hcbe1;
aud[7927]=16'hcbd5;
aud[7928]=16'hcbc9;
aud[7929]=16'hcbbc;
aud[7930]=16'hcbb0;
aud[7931]=16'hcba3;
aud[7932]=16'hcb97;
aud[7933]=16'hcb8b;
aud[7934]=16'hcb7f;
aud[7935]=16'hcb72;
aud[7936]=16'hcb66;
aud[7937]=16'hcb5a;
aud[7938]=16'hcb4e;
aud[7939]=16'hcb42;
aud[7940]=16'hcb35;
aud[7941]=16'hcb29;
aud[7942]=16'hcb1d;
aud[7943]=16'hcb11;
aud[7944]=16'hcb05;
aud[7945]=16'hcaf9;
aud[7946]=16'hcaed;
aud[7947]=16'hcae1;
aud[7948]=16'hcad5;
aud[7949]=16'hcac9;
aud[7950]=16'hcabd;
aud[7951]=16'hcab1;
aud[7952]=16'hcaa6;
aud[7953]=16'hca9a;
aud[7954]=16'hca8e;
aud[7955]=16'hca82;
aud[7956]=16'hca76;
aud[7957]=16'hca6b;
aud[7958]=16'hca5f;
aud[7959]=16'hca53;
aud[7960]=16'hca48;
aud[7961]=16'hca3c;
aud[7962]=16'hca30;
aud[7963]=16'hca25;
aud[7964]=16'hca19;
aud[7965]=16'hca0e;
aud[7966]=16'hca02;
aud[7967]=16'hc9f7;
aud[7968]=16'hc9eb;
aud[7969]=16'hc9e0;
aud[7970]=16'hc9d4;
aud[7971]=16'hc9c9;
aud[7972]=16'hc9bd;
aud[7973]=16'hc9b2;
aud[7974]=16'hc9a7;
aud[7975]=16'hc99b;
aud[7976]=16'hc990;
aud[7977]=16'hc985;
aud[7978]=16'hc97a;
aud[7979]=16'hc96e;
aud[7980]=16'hc963;
aud[7981]=16'hc958;
aud[7982]=16'hc94d;
aud[7983]=16'hc942;
aud[7984]=16'hc937;
aud[7985]=16'hc92c;
aud[7986]=16'hc920;
aud[7987]=16'hc915;
aud[7988]=16'hc90a;
aud[7989]=16'hc8ff;
aud[7990]=16'hc8f5;
aud[7991]=16'hc8ea;
aud[7992]=16'hc8df;
aud[7993]=16'hc8d4;
aud[7994]=16'hc8c9;
aud[7995]=16'hc8be;
aud[7996]=16'hc8b3;
aud[7997]=16'hc8a9;
aud[7998]=16'hc89e;
aud[7999]=16'hc893;
aud[8000]=16'hc888;
aud[8001]=16'hc87e;
aud[8002]=16'hc873;
aud[8003]=16'hc868;
aud[8004]=16'hc85e;
aud[8005]=16'hc853;
aud[8006]=16'hc849;
aud[8007]=16'hc83e;
aud[8008]=16'hc834;
aud[8009]=16'hc829;
aud[8010]=16'hc81f;
aud[8011]=16'hc814;
aud[8012]=16'hc80a;
aud[8013]=16'hc7ff;
aud[8014]=16'hc7f5;
aud[8015]=16'hc7eb;
aud[8016]=16'hc7e0;
aud[8017]=16'hc7d6;
aud[8018]=16'hc7cc;
aud[8019]=16'hc7c1;
aud[8020]=16'hc7b7;
aud[8021]=16'hc7ad;
aud[8022]=16'hc7a3;
aud[8023]=16'hc799;
aud[8024]=16'hc78f;
aud[8025]=16'hc785;
aud[8026]=16'hc77a;
aud[8027]=16'hc770;
aud[8028]=16'hc766;
aud[8029]=16'hc75c;
aud[8030]=16'hc752;
aud[8031]=16'hc748;
aud[8032]=16'hc73f;
aud[8033]=16'hc735;
aud[8034]=16'hc72b;
aud[8035]=16'hc721;
aud[8036]=16'hc717;
aud[8037]=16'hc70d;
aud[8038]=16'hc703;
aud[8039]=16'hc6fa;
aud[8040]=16'hc6f0;
aud[8041]=16'hc6e6;
aud[8042]=16'hc6dd;
aud[8043]=16'hc6d3;
aud[8044]=16'hc6c9;
aud[8045]=16'hc6c0;
aud[8046]=16'hc6b6;
aud[8047]=16'hc6ad;
aud[8048]=16'hc6a3;
aud[8049]=16'hc69a;
aud[8050]=16'hc690;
aud[8051]=16'hc687;
aud[8052]=16'hc67d;
aud[8053]=16'hc674;
aud[8054]=16'hc66b;
aud[8055]=16'hc661;
aud[8056]=16'hc658;
aud[8057]=16'hc64f;
aud[8058]=16'hc645;
aud[8059]=16'hc63c;
aud[8060]=16'hc633;
aud[8061]=16'hc62a;
aud[8062]=16'hc620;
aud[8063]=16'hc617;
aud[8064]=16'hc60e;
aud[8065]=16'hc605;
aud[8066]=16'hc5fc;
aud[8067]=16'hc5f3;
aud[8068]=16'hc5ea;
aud[8069]=16'hc5e1;
aud[8070]=16'hc5d8;
aud[8071]=16'hc5cf;
aud[8072]=16'hc5c6;
aud[8073]=16'hc5bd;
aud[8074]=16'hc5b4;
aud[8075]=16'hc5ac;
aud[8076]=16'hc5a3;
aud[8077]=16'hc59a;
aud[8078]=16'hc591;
aud[8079]=16'hc588;
aud[8080]=16'hc580;
aud[8081]=16'hc577;
aud[8082]=16'hc56e;
aud[8083]=16'hc566;
aud[8084]=16'hc55d;
aud[8085]=16'hc555;
aud[8086]=16'hc54c;
aud[8087]=16'hc544;
aud[8088]=16'hc53b;
aud[8089]=16'hc533;
aud[8090]=16'hc52a;
aud[8091]=16'hc522;
aud[8092]=16'hc519;
aud[8093]=16'hc511;
aud[8094]=16'hc509;
aud[8095]=16'hc500;
aud[8096]=16'hc4f8;
aud[8097]=16'hc4f0;
aud[8098]=16'hc4e7;
aud[8099]=16'hc4df;
aud[8100]=16'hc4d7;
aud[8101]=16'hc4cf;
aud[8102]=16'hc4c7;
aud[8103]=16'hc4bf;
aud[8104]=16'hc4b6;
aud[8105]=16'hc4ae;
aud[8106]=16'hc4a6;
aud[8107]=16'hc49e;
aud[8108]=16'hc496;
aud[8109]=16'hc48e;
aud[8110]=16'hc486;
aud[8111]=16'hc47f;
aud[8112]=16'hc477;
aud[8113]=16'hc46f;
aud[8114]=16'hc467;
aud[8115]=16'hc45f;
aud[8116]=16'hc457;
aud[8117]=16'hc450;
aud[8118]=16'hc448;
aud[8119]=16'hc440;
aud[8120]=16'hc439;
aud[8121]=16'hc431;
aud[8122]=16'hc429;
aud[8123]=16'hc422;
aud[8124]=16'hc41a;
aud[8125]=16'hc413;
aud[8126]=16'hc40b;
aud[8127]=16'hc404;
aud[8128]=16'hc3fc;
aud[8129]=16'hc3f5;
aud[8130]=16'hc3ed;
aud[8131]=16'hc3e6;
aud[8132]=16'hc3df;
aud[8133]=16'hc3d7;
aud[8134]=16'hc3d0;
aud[8135]=16'hc3c9;
aud[8136]=16'hc3c1;
aud[8137]=16'hc3ba;
aud[8138]=16'hc3b3;
aud[8139]=16'hc3ac;
aud[8140]=16'hc3a5;
aud[8141]=16'hc39d;
aud[8142]=16'hc396;
aud[8143]=16'hc38f;
aud[8144]=16'hc388;
aud[8145]=16'hc381;
aud[8146]=16'hc37a;
aud[8147]=16'hc373;
aud[8148]=16'hc36c;
aud[8149]=16'hc365;
aud[8150]=16'hc35f;
aud[8151]=16'hc358;
aud[8152]=16'hc351;
aud[8153]=16'hc34a;
aud[8154]=16'hc343;
aud[8155]=16'hc33d;
aud[8156]=16'hc336;
aud[8157]=16'hc32f;
aud[8158]=16'hc329;
aud[8159]=16'hc322;
aud[8160]=16'hc31b;
aud[8161]=16'hc315;
aud[8162]=16'hc30e;
aud[8163]=16'hc308;
aud[8164]=16'hc301;
aud[8165]=16'hc2fb;
aud[8166]=16'hc2f4;
aud[8167]=16'hc2ee;
aud[8168]=16'hc2e7;
aud[8169]=16'hc2e1;
aud[8170]=16'hc2db;
aud[8171]=16'hc2d4;
aud[8172]=16'hc2ce;
aud[8173]=16'hc2c8;
aud[8174]=16'hc2c1;
aud[8175]=16'hc2bb;
aud[8176]=16'hc2b5;
aud[8177]=16'hc2af;
aud[8178]=16'hc2a9;
aud[8179]=16'hc2a3;
aud[8180]=16'hc29d;
aud[8181]=16'hc297;
aud[8182]=16'hc291;
aud[8183]=16'hc28b;
aud[8184]=16'hc285;
aud[8185]=16'hc27f;
aud[8186]=16'hc279;
aud[8187]=16'hc273;
aud[8188]=16'hc26d;
aud[8189]=16'hc267;
aud[8190]=16'hc261;
aud[8191]=16'hc25c;
aud[8192]=16'hc256;
aud[8193]=16'hc250;
aud[8194]=16'hc24a;
aud[8195]=16'hc245;
aud[8196]=16'hc23f;
aud[8197]=16'hc239;
aud[8198]=16'hc234;
aud[8199]=16'hc22e;
aud[8200]=16'hc229;
aud[8201]=16'hc223;
aud[8202]=16'hc21e;
aud[8203]=16'hc218;
aud[8204]=16'hc213;
aud[8205]=16'hc20d;
aud[8206]=16'hc208;
aud[8207]=16'hc203;
aud[8208]=16'hc1fd;
aud[8209]=16'hc1f8;
aud[8210]=16'hc1f3;
aud[8211]=16'hc1ee;
aud[8212]=16'hc1e8;
aud[8213]=16'hc1e3;
aud[8214]=16'hc1de;
aud[8215]=16'hc1d9;
aud[8216]=16'hc1d4;
aud[8217]=16'hc1cf;
aud[8218]=16'hc1ca;
aud[8219]=16'hc1c5;
aud[8220]=16'hc1c0;
aud[8221]=16'hc1bb;
aud[8222]=16'hc1b6;
aud[8223]=16'hc1b1;
aud[8224]=16'hc1ac;
aud[8225]=16'hc1a7;
aud[8226]=16'hc1a2;
aud[8227]=16'hc19e;
aud[8228]=16'hc199;
aud[8229]=16'hc194;
aud[8230]=16'hc18f;
aud[8231]=16'hc18b;
aud[8232]=16'hc186;
aud[8233]=16'hc181;
aud[8234]=16'hc17d;
aud[8235]=16'hc178;
aud[8236]=16'hc174;
aud[8237]=16'hc16f;
aud[8238]=16'hc16b;
aud[8239]=16'hc166;
aud[8240]=16'hc162;
aud[8241]=16'hc15d;
aud[8242]=16'hc159;
aud[8243]=16'hc154;
aud[8244]=16'hc150;
aud[8245]=16'hc14c;
aud[8246]=16'hc147;
aud[8247]=16'hc143;
aud[8248]=16'hc13f;
aud[8249]=16'hc13b;
aud[8250]=16'hc137;
aud[8251]=16'hc133;
aud[8252]=16'hc12e;
aud[8253]=16'hc12a;
aud[8254]=16'hc126;
aud[8255]=16'hc122;
aud[8256]=16'hc11e;
aud[8257]=16'hc11a;
aud[8258]=16'hc116;
aud[8259]=16'hc112;
aud[8260]=16'hc10e;
aud[8261]=16'hc10b;
aud[8262]=16'hc107;
aud[8263]=16'hc103;
aud[8264]=16'hc0ff;
aud[8265]=16'hc0fb;
aud[8266]=16'hc0f8;
aud[8267]=16'hc0f4;
aud[8268]=16'hc0f0;
aud[8269]=16'hc0ed;
aud[8270]=16'hc0e9;
aud[8271]=16'hc0e5;
aud[8272]=16'hc0e2;
aud[8273]=16'hc0de;
aud[8274]=16'hc0db;
aud[8275]=16'hc0d7;
aud[8276]=16'hc0d4;
aud[8277]=16'hc0d0;
aud[8278]=16'hc0cd;
aud[8279]=16'hc0ca;
aud[8280]=16'hc0c6;
aud[8281]=16'hc0c3;
aud[8282]=16'hc0c0;
aud[8283]=16'hc0bd;
aud[8284]=16'hc0b9;
aud[8285]=16'hc0b6;
aud[8286]=16'hc0b3;
aud[8287]=16'hc0b0;
aud[8288]=16'hc0ad;
aud[8289]=16'hc0aa;
aud[8290]=16'hc0a6;
aud[8291]=16'hc0a3;
aud[8292]=16'hc0a0;
aud[8293]=16'hc09d;
aud[8294]=16'hc09b;
aud[8295]=16'hc098;
aud[8296]=16'hc095;
aud[8297]=16'hc092;
aud[8298]=16'hc08f;
aud[8299]=16'hc08c;
aud[8300]=16'hc089;
aud[8301]=16'hc087;
aud[8302]=16'hc084;
aud[8303]=16'hc081;
aud[8304]=16'hc07f;
aud[8305]=16'hc07c;
aud[8306]=16'hc079;
aud[8307]=16'hc077;
aud[8308]=16'hc074;
aud[8309]=16'hc072;
aud[8310]=16'hc06f;
aud[8311]=16'hc06d;
aud[8312]=16'hc06a;
aud[8313]=16'hc068;
aud[8314]=16'hc065;
aud[8315]=16'hc063;
aud[8316]=16'hc061;
aud[8317]=16'hc05e;
aud[8318]=16'hc05c;
aud[8319]=16'hc05a;
aud[8320]=16'hc058;
aud[8321]=16'hc055;
aud[8322]=16'hc053;
aud[8323]=16'hc051;
aud[8324]=16'hc04f;
aud[8325]=16'hc04d;
aud[8326]=16'hc04b;
aud[8327]=16'hc049;
aud[8328]=16'hc047;
aud[8329]=16'hc045;
aud[8330]=16'hc043;
aud[8331]=16'hc041;
aud[8332]=16'hc03f;
aud[8333]=16'hc03d;
aud[8334]=16'hc03b;
aud[8335]=16'hc039;
aud[8336]=16'hc038;
aud[8337]=16'hc036;
aud[8338]=16'hc034;
aud[8339]=16'hc033;
aud[8340]=16'hc031;
aud[8341]=16'hc02f;
aud[8342]=16'hc02e;
aud[8343]=16'hc02c;
aud[8344]=16'hc02a;
aud[8345]=16'hc029;
aud[8346]=16'hc027;
aud[8347]=16'hc026;
aud[8348]=16'hc024;
aud[8349]=16'hc023;
aud[8350]=16'hc022;
aud[8351]=16'hc020;
aud[8352]=16'hc01f;
aud[8353]=16'hc01e;
aud[8354]=16'hc01c;
aud[8355]=16'hc01b;
aud[8356]=16'hc01a;
aud[8357]=16'hc019;
aud[8358]=16'hc018;
aud[8359]=16'hc016;
aud[8360]=16'hc015;
aud[8361]=16'hc014;
aud[8362]=16'hc013;
aud[8363]=16'hc012;
aud[8364]=16'hc011;
aud[8365]=16'hc010;
aud[8366]=16'hc00f;
aud[8367]=16'hc00e;
aud[8368]=16'hc00d;
aud[8369]=16'hc00d;
aud[8370]=16'hc00c;
aud[8371]=16'hc00b;
aud[8372]=16'hc00a;
aud[8373]=16'hc009;
aud[8374]=16'hc009;
aud[8375]=16'hc008;
aud[8376]=16'hc007;
aud[8377]=16'hc007;
aud[8378]=16'hc006;
aud[8379]=16'hc006;
aud[8380]=16'hc005;
aud[8381]=16'hc005;
aud[8382]=16'hc004;
aud[8383]=16'hc004;
aud[8384]=16'hc003;
aud[8385]=16'hc003;
aud[8386]=16'hc002;
aud[8387]=16'hc002;
aud[8388]=16'hc002;
aud[8389]=16'hc001;
aud[8390]=16'hc001;
aud[8391]=16'hc001;
aud[8392]=16'hc001;
aud[8393]=16'hc001;
aud[8394]=16'hc000;
aud[8395]=16'hc000;
aud[8396]=16'hc000;
aud[8397]=16'hc000;
aud[8398]=16'hc000;
aud[8399]=16'hc000;
aud[8400]=16'hc000;
aud[8401]=16'hc000;
aud[8402]=16'hc000;
aud[8403]=16'hc000;
aud[8404]=16'hc000;
aud[8405]=16'hc001;
aud[8406]=16'hc001;
aud[8407]=16'hc001;
aud[8408]=16'hc001;
aud[8409]=16'hc001;
aud[8410]=16'hc002;
aud[8411]=16'hc002;
aud[8412]=16'hc002;
aud[8413]=16'hc003;
aud[8414]=16'hc003;
aud[8415]=16'hc004;
aud[8416]=16'hc004;
aud[8417]=16'hc005;
aud[8418]=16'hc005;
aud[8419]=16'hc006;
aud[8420]=16'hc006;
aud[8421]=16'hc007;
aud[8422]=16'hc007;
aud[8423]=16'hc008;
aud[8424]=16'hc009;
aud[8425]=16'hc009;
aud[8426]=16'hc00a;
aud[8427]=16'hc00b;
aud[8428]=16'hc00c;
aud[8429]=16'hc00d;
aud[8430]=16'hc00d;
aud[8431]=16'hc00e;
aud[8432]=16'hc00f;
aud[8433]=16'hc010;
aud[8434]=16'hc011;
aud[8435]=16'hc012;
aud[8436]=16'hc013;
aud[8437]=16'hc014;
aud[8438]=16'hc015;
aud[8439]=16'hc016;
aud[8440]=16'hc018;
aud[8441]=16'hc019;
aud[8442]=16'hc01a;
aud[8443]=16'hc01b;
aud[8444]=16'hc01c;
aud[8445]=16'hc01e;
aud[8446]=16'hc01f;
aud[8447]=16'hc020;
aud[8448]=16'hc022;
aud[8449]=16'hc023;
aud[8450]=16'hc024;
aud[8451]=16'hc026;
aud[8452]=16'hc027;
aud[8453]=16'hc029;
aud[8454]=16'hc02a;
aud[8455]=16'hc02c;
aud[8456]=16'hc02e;
aud[8457]=16'hc02f;
aud[8458]=16'hc031;
aud[8459]=16'hc033;
aud[8460]=16'hc034;
aud[8461]=16'hc036;
aud[8462]=16'hc038;
aud[8463]=16'hc039;
aud[8464]=16'hc03b;
aud[8465]=16'hc03d;
aud[8466]=16'hc03f;
aud[8467]=16'hc041;
aud[8468]=16'hc043;
aud[8469]=16'hc045;
aud[8470]=16'hc047;
aud[8471]=16'hc049;
aud[8472]=16'hc04b;
aud[8473]=16'hc04d;
aud[8474]=16'hc04f;
aud[8475]=16'hc051;
aud[8476]=16'hc053;
aud[8477]=16'hc055;
aud[8478]=16'hc058;
aud[8479]=16'hc05a;
aud[8480]=16'hc05c;
aud[8481]=16'hc05e;
aud[8482]=16'hc061;
aud[8483]=16'hc063;
aud[8484]=16'hc065;
aud[8485]=16'hc068;
aud[8486]=16'hc06a;
aud[8487]=16'hc06d;
aud[8488]=16'hc06f;
aud[8489]=16'hc072;
aud[8490]=16'hc074;
aud[8491]=16'hc077;
aud[8492]=16'hc079;
aud[8493]=16'hc07c;
aud[8494]=16'hc07f;
aud[8495]=16'hc081;
aud[8496]=16'hc084;
aud[8497]=16'hc087;
aud[8498]=16'hc089;
aud[8499]=16'hc08c;
aud[8500]=16'hc08f;
aud[8501]=16'hc092;
aud[8502]=16'hc095;
aud[8503]=16'hc098;
aud[8504]=16'hc09b;
aud[8505]=16'hc09d;
aud[8506]=16'hc0a0;
aud[8507]=16'hc0a3;
aud[8508]=16'hc0a6;
aud[8509]=16'hc0aa;
aud[8510]=16'hc0ad;
aud[8511]=16'hc0b0;
aud[8512]=16'hc0b3;
aud[8513]=16'hc0b6;
aud[8514]=16'hc0b9;
aud[8515]=16'hc0bd;
aud[8516]=16'hc0c0;
aud[8517]=16'hc0c3;
aud[8518]=16'hc0c6;
aud[8519]=16'hc0ca;
aud[8520]=16'hc0cd;
aud[8521]=16'hc0d0;
aud[8522]=16'hc0d4;
aud[8523]=16'hc0d7;
aud[8524]=16'hc0db;
aud[8525]=16'hc0de;
aud[8526]=16'hc0e2;
aud[8527]=16'hc0e5;
aud[8528]=16'hc0e9;
aud[8529]=16'hc0ed;
aud[8530]=16'hc0f0;
aud[8531]=16'hc0f4;
aud[8532]=16'hc0f8;
aud[8533]=16'hc0fb;
aud[8534]=16'hc0ff;
aud[8535]=16'hc103;
aud[8536]=16'hc107;
aud[8537]=16'hc10b;
aud[8538]=16'hc10e;
aud[8539]=16'hc112;
aud[8540]=16'hc116;
aud[8541]=16'hc11a;
aud[8542]=16'hc11e;
aud[8543]=16'hc122;
aud[8544]=16'hc126;
aud[8545]=16'hc12a;
aud[8546]=16'hc12e;
aud[8547]=16'hc133;
aud[8548]=16'hc137;
aud[8549]=16'hc13b;
aud[8550]=16'hc13f;
aud[8551]=16'hc143;
aud[8552]=16'hc147;
aud[8553]=16'hc14c;
aud[8554]=16'hc150;
aud[8555]=16'hc154;
aud[8556]=16'hc159;
aud[8557]=16'hc15d;
aud[8558]=16'hc162;
aud[8559]=16'hc166;
aud[8560]=16'hc16b;
aud[8561]=16'hc16f;
aud[8562]=16'hc174;
aud[8563]=16'hc178;
aud[8564]=16'hc17d;
aud[8565]=16'hc181;
aud[8566]=16'hc186;
aud[8567]=16'hc18b;
aud[8568]=16'hc18f;
aud[8569]=16'hc194;
aud[8570]=16'hc199;
aud[8571]=16'hc19e;
aud[8572]=16'hc1a2;
aud[8573]=16'hc1a7;
aud[8574]=16'hc1ac;
aud[8575]=16'hc1b1;
aud[8576]=16'hc1b6;
aud[8577]=16'hc1bb;
aud[8578]=16'hc1c0;
aud[8579]=16'hc1c5;
aud[8580]=16'hc1ca;
aud[8581]=16'hc1cf;
aud[8582]=16'hc1d4;
aud[8583]=16'hc1d9;
aud[8584]=16'hc1de;
aud[8585]=16'hc1e3;
aud[8586]=16'hc1e8;
aud[8587]=16'hc1ee;
aud[8588]=16'hc1f3;
aud[8589]=16'hc1f8;
aud[8590]=16'hc1fd;
aud[8591]=16'hc203;
aud[8592]=16'hc208;
aud[8593]=16'hc20d;
aud[8594]=16'hc213;
aud[8595]=16'hc218;
aud[8596]=16'hc21e;
aud[8597]=16'hc223;
aud[8598]=16'hc229;
aud[8599]=16'hc22e;
aud[8600]=16'hc234;
aud[8601]=16'hc239;
aud[8602]=16'hc23f;
aud[8603]=16'hc245;
aud[8604]=16'hc24a;
aud[8605]=16'hc250;
aud[8606]=16'hc256;
aud[8607]=16'hc25c;
aud[8608]=16'hc261;
aud[8609]=16'hc267;
aud[8610]=16'hc26d;
aud[8611]=16'hc273;
aud[8612]=16'hc279;
aud[8613]=16'hc27f;
aud[8614]=16'hc285;
aud[8615]=16'hc28b;
aud[8616]=16'hc291;
aud[8617]=16'hc297;
aud[8618]=16'hc29d;
aud[8619]=16'hc2a3;
aud[8620]=16'hc2a9;
aud[8621]=16'hc2af;
aud[8622]=16'hc2b5;
aud[8623]=16'hc2bb;
aud[8624]=16'hc2c1;
aud[8625]=16'hc2c8;
aud[8626]=16'hc2ce;
aud[8627]=16'hc2d4;
aud[8628]=16'hc2db;
aud[8629]=16'hc2e1;
aud[8630]=16'hc2e7;
aud[8631]=16'hc2ee;
aud[8632]=16'hc2f4;
aud[8633]=16'hc2fb;
aud[8634]=16'hc301;
aud[8635]=16'hc308;
aud[8636]=16'hc30e;
aud[8637]=16'hc315;
aud[8638]=16'hc31b;
aud[8639]=16'hc322;
aud[8640]=16'hc329;
aud[8641]=16'hc32f;
aud[8642]=16'hc336;
aud[8643]=16'hc33d;
aud[8644]=16'hc343;
aud[8645]=16'hc34a;
aud[8646]=16'hc351;
aud[8647]=16'hc358;
aud[8648]=16'hc35f;
aud[8649]=16'hc365;
aud[8650]=16'hc36c;
aud[8651]=16'hc373;
aud[8652]=16'hc37a;
aud[8653]=16'hc381;
aud[8654]=16'hc388;
aud[8655]=16'hc38f;
aud[8656]=16'hc396;
aud[8657]=16'hc39d;
aud[8658]=16'hc3a5;
aud[8659]=16'hc3ac;
aud[8660]=16'hc3b3;
aud[8661]=16'hc3ba;
aud[8662]=16'hc3c1;
aud[8663]=16'hc3c9;
aud[8664]=16'hc3d0;
aud[8665]=16'hc3d7;
aud[8666]=16'hc3df;
aud[8667]=16'hc3e6;
aud[8668]=16'hc3ed;
aud[8669]=16'hc3f5;
aud[8670]=16'hc3fc;
aud[8671]=16'hc404;
aud[8672]=16'hc40b;
aud[8673]=16'hc413;
aud[8674]=16'hc41a;
aud[8675]=16'hc422;
aud[8676]=16'hc429;
aud[8677]=16'hc431;
aud[8678]=16'hc439;
aud[8679]=16'hc440;
aud[8680]=16'hc448;
aud[8681]=16'hc450;
aud[8682]=16'hc457;
aud[8683]=16'hc45f;
aud[8684]=16'hc467;
aud[8685]=16'hc46f;
aud[8686]=16'hc477;
aud[8687]=16'hc47f;
aud[8688]=16'hc486;
aud[8689]=16'hc48e;
aud[8690]=16'hc496;
aud[8691]=16'hc49e;
aud[8692]=16'hc4a6;
aud[8693]=16'hc4ae;
aud[8694]=16'hc4b6;
aud[8695]=16'hc4bf;
aud[8696]=16'hc4c7;
aud[8697]=16'hc4cf;
aud[8698]=16'hc4d7;
aud[8699]=16'hc4df;
aud[8700]=16'hc4e7;
aud[8701]=16'hc4f0;
aud[8702]=16'hc4f8;
aud[8703]=16'hc500;
aud[8704]=16'hc509;
aud[8705]=16'hc511;
aud[8706]=16'hc519;
aud[8707]=16'hc522;
aud[8708]=16'hc52a;
aud[8709]=16'hc533;
aud[8710]=16'hc53b;
aud[8711]=16'hc544;
aud[8712]=16'hc54c;
aud[8713]=16'hc555;
aud[8714]=16'hc55d;
aud[8715]=16'hc566;
aud[8716]=16'hc56e;
aud[8717]=16'hc577;
aud[8718]=16'hc580;
aud[8719]=16'hc588;
aud[8720]=16'hc591;
aud[8721]=16'hc59a;
aud[8722]=16'hc5a3;
aud[8723]=16'hc5ac;
aud[8724]=16'hc5b4;
aud[8725]=16'hc5bd;
aud[8726]=16'hc5c6;
aud[8727]=16'hc5cf;
aud[8728]=16'hc5d8;
aud[8729]=16'hc5e1;
aud[8730]=16'hc5ea;
aud[8731]=16'hc5f3;
aud[8732]=16'hc5fc;
aud[8733]=16'hc605;
aud[8734]=16'hc60e;
aud[8735]=16'hc617;
aud[8736]=16'hc620;
aud[8737]=16'hc62a;
aud[8738]=16'hc633;
aud[8739]=16'hc63c;
aud[8740]=16'hc645;
aud[8741]=16'hc64f;
aud[8742]=16'hc658;
aud[8743]=16'hc661;
aud[8744]=16'hc66b;
aud[8745]=16'hc674;
aud[8746]=16'hc67d;
aud[8747]=16'hc687;
aud[8748]=16'hc690;
aud[8749]=16'hc69a;
aud[8750]=16'hc6a3;
aud[8751]=16'hc6ad;
aud[8752]=16'hc6b6;
aud[8753]=16'hc6c0;
aud[8754]=16'hc6c9;
aud[8755]=16'hc6d3;
aud[8756]=16'hc6dd;
aud[8757]=16'hc6e6;
aud[8758]=16'hc6f0;
aud[8759]=16'hc6fa;
aud[8760]=16'hc703;
aud[8761]=16'hc70d;
aud[8762]=16'hc717;
aud[8763]=16'hc721;
aud[8764]=16'hc72b;
aud[8765]=16'hc735;
aud[8766]=16'hc73f;
aud[8767]=16'hc748;
aud[8768]=16'hc752;
aud[8769]=16'hc75c;
aud[8770]=16'hc766;
aud[8771]=16'hc770;
aud[8772]=16'hc77a;
aud[8773]=16'hc785;
aud[8774]=16'hc78f;
aud[8775]=16'hc799;
aud[8776]=16'hc7a3;
aud[8777]=16'hc7ad;
aud[8778]=16'hc7b7;
aud[8779]=16'hc7c1;
aud[8780]=16'hc7cc;
aud[8781]=16'hc7d6;
aud[8782]=16'hc7e0;
aud[8783]=16'hc7eb;
aud[8784]=16'hc7f5;
aud[8785]=16'hc7ff;
aud[8786]=16'hc80a;
aud[8787]=16'hc814;
aud[8788]=16'hc81f;
aud[8789]=16'hc829;
aud[8790]=16'hc834;
aud[8791]=16'hc83e;
aud[8792]=16'hc849;
aud[8793]=16'hc853;
aud[8794]=16'hc85e;
aud[8795]=16'hc868;
aud[8796]=16'hc873;
aud[8797]=16'hc87e;
aud[8798]=16'hc888;
aud[8799]=16'hc893;
aud[8800]=16'hc89e;
aud[8801]=16'hc8a9;
aud[8802]=16'hc8b3;
aud[8803]=16'hc8be;
aud[8804]=16'hc8c9;
aud[8805]=16'hc8d4;
aud[8806]=16'hc8df;
aud[8807]=16'hc8ea;
aud[8808]=16'hc8f5;
aud[8809]=16'hc8ff;
aud[8810]=16'hc90a;
aud[8811]=16'hc915;
aud[8812]=16'hc920;
aud[8813]=16'hc92c;
aud[8814]=16'hc937;
aud[8815]=16'hc942;
aud[8816]=16'hc94d;
aud[8817]=16'hc958;
aud[8818]=16'hc963;
aud[8819]=16'hc96e;
aud[8820]=16'hc97a;
aud[8821]=16'hc985;
aud[8822]=16'hc990;
aud[8823]=16'hc99b;
aud[8824]=16'hc9a7;
aud[8825]=16'hc9b2;
aud[8826]=16'hc9bd;
aud[8827]=16'hc9c9;
aud[8828]=16'hc9d4;
aud[8829]=16'hc9e0;
aud[8830]=16'hc9eb;
aud[8831]=16'hc9f7;
aud[8832]=16'hca02;
aud[8833]=16'hca0e;
aud[8834]=16'hca19;
aud[8835]=16'hca25;
aud[8836]=16'hca30;
aud[8837]=16'hca3c;
aud[8838]=16'hca48;
aud[8839]=16'hca53;
aud[8840]=16'hca5f;
aud[8841]=16'hca6b;
aud[8842]=16'hca76;
aud[8843]=16'hca82;
aud[8844]=16'hca8e;
aud[8845]=16'hca9a;
aud[8846]=16'hcaa6;
aud[8847]=16'hcab1;
aud[8848]=16'hcabd;
aud[8849]=16'hcac9;
aud[8850]=16'hcad5;
aud[8851]=16'hcae1;
aud[8852]=16'hcaed;
aud[8853]=16'hcaf9;
aud[8854]=16'hcb05;
aud[8855]=16'hcb11;
aud[8856]=16'hcb1d;
aud[8857]=16'hcb29;
aud[8858]=16'hcb35;
aud[8859]=16'hcb42;
aud[8860]=16'hcb4e;
aud[8861]=16'hcb5a;
aud[8862]=16'hcb66;
aud[8863]=16'hcb72;
aud[8864]=16'hcb7f;
aud[8865]=16'hcb8b;
aud[8866]=16'hcb97;
aud[8867]=16'hcba3;
aud[8868]=16'hcbb0;
aud[8869]=16'hcbbc;
aud[8870]=16'hcbc9;
aud[8871]=16'hcbd5;
aud[8872]=16'hcbe1;
aud[8873]=16'hcbee;
aud[8874]=16'hcbfa;
aud[8875]=16'hcc07;
aud[8876]=16'hcc13;
aud[8877]=16'hcc20;
aud[8878]=16'hcc2c;
aud[8879]=16'hcc39;
aud[8880]=16'hcc46;
aud[8881]=16'hcc52;
aud[8882]=16'hcc5f;
aud[8883]=16'hcc6c;
aud[8884]=16'hcc78;
aud[8885]=16'hcc85;
aud[8886]=16'hcc92;
aud[8887]=16'hcc9f;
aud[8888]=16'hccab;
aud[8889]=16'hccb8;
aud[8890]=16'hccc5;
aud[8891]=16'hccd2;
aud[8892]=16'hccdf;
aud[8893]=16'hccec;
aud[8894]=16'hccf9;
aud[8895]=16'hcd06;
aud[8896]=16'hcd13;
aud[8897]=16'hcd20;
aud[8898]=16'hcd2d;
aud[8899]=16'hcd3a;
aud[8900]=16'hcd47;
aud[8901]=16'hcd54;
aud[8902]=16'hcd61;
aud[8903]=16'hcd6e;
aud[8904]=16'hcd7b;
aud[8905]=16'hcd88;
aud[8906]=16'hcd96;
aud[8907]=16'hcda3;
aud[8908]=16'hcdb0;
aud[8909]=16'hcdbd;
aud[8910]=16'hcdcb;
aud[8911]=16'hcdd8;
aud[8912]=16'hcde5;
aud[8913]=16'hcdf3;
aud[8914]=16'hce00;
aud[8915]=16'hce0d;
aud[8916]=16'hce1b;
aud[8917]=16'hce28;
aud[8918]=16'hce36;
aud[8919]=16'hce43;
aud[8920]=16'hce51;
aud[8921]=16'hce5e;
aud[8922]=16'hce6c;
aud[8923]=16'hce79;
aud[8924]=16'hce87;
aud[8925]=16'hce95;
aud[8926]=16'hcea2;
aud[8927]=16'hceb0;
aud[8928]=16'hcebe;
aud[8929]=16'hcecb;
aud[8930]=16'hced9;
aud[8931]=16'hcee7;
aud[8932]=16'hcef5;
aud[8933]=16'hcf02;
aud[8934]=16'hcf10;
aud[8935]=16'hcf1e;
aud[8936]=16'hcf2c;
aud[8937]=16'hcf3a;
aud[8938]=16'hcf48;
aud[8939]=16'hcf56;
aud[8940]=16'hcf63;
aud[8941]=16'hcf71;
aud[8942]=16'hcf7f;
aud[8943]=16'hcf8d;
aud[8944]=16'hcf9b;
aud[8945]=16'hcfa9;
aud[8946]=16'hcfb8;
aud[8947]=16'hcfc6;
aud[8948]=16'hcfd4;
aud[8949]=16'hcfe2;
aud[8950]=16'hcff0;
aud[8951]=16'hcffe;
aud[8952]=16'hd00c;
aud[8953]=16'hd01b;
aud[8954]=16'hd029;
aud[8955]=16'hd037;
aud[8956]=16'hd045;
aud[8957]=16'hd054;
aud[8958]=16'hd062;
aud[8959]=16'hd070;
aud[8960]=16'hd07f;
aud[8961]=16'hd08d;
aud[8962]=16'hd09b;
aud[8963]=16'hd0aa;
aud[8964]=16'hd0b8;
aud[8965]=16'hd0c7;
aud[8966]=16'hd0d5;
aud[8967]=16'hd0e4;
aud[8968]=16'hd0f2;
aud[8969]=16'hd101;
aud[8970]=16'hd10f;
aud[8971]=16'hd11e;
aud[8972]=16'hd12d;
aud[8973]=16'hd13b;
aud[8974]=16'hd14a;
aud[8975]=16'hd159;
aud[8976]=16'hd167;
aud[8977]=16'hd176;
aud[8978]=16'hd185;
aud[8979]=16'hd193;
aud[8980]=16'hd1a2;
aud[8981]=16'hd1b1;
aud[8982]=16'hd1c0;
aud[8983]=16'hd1cf;
aud[8984]=16'hd1de;
aud[8985]=16'hd1ec;
aud[8986]=16'hd1fb;
aud[8987]=16'hd20a;
aud[8988]=16'hd219;
aud[8989]=16'hd228;
aud[8990]=16'hd237;
aud[8991]=16'hd246;
aud[8992]=16'hd255;
aud[8993]=16'hd264;
aud[8994]=16'hd273;
aud[8995]=16'hd282;
aud[8996]=16'hd291;
aud[8997]=16'hd2a0;
aud[8998]=16'hd2b0;
aud[8999]=16'hd2bf;
aud[9000]=16'hd2ce;
aud[9001]=16'hd2dd;
aud[9002]=16'hd2ec;
aud[9003]=16'hd2fc;
aud[9004]=16'hd30b;
aud[9005]=16'hd31a;
aud[9006]=16'hd329;
aud[9007]=16'hd339;
aud[9008]=16'hd348;
aud[9009]=16'hd357;
aud[9010]=16'hd367;
aud[9011]=16'hd376;
aud[9012]=16'hd386;
aud[9013]=16'hd395;
aud[9014]=16'hd3a4;
aud[9015]=16'hd3b4;
aud[9016]=16'hd3c3;
aud[9017]=16'hd3d3;
aud[9018]=16'hd3e2;
aud[9019]=16'hd3f2;
aud[9020]=16'hd402;
aud[9021]=16'hd411;
aud[9022]=16'hd421;
aud[9023]=16'hd430;
aud[9024]=16'hd440;
aud[9025]=16'hd450;
aud[9026]=16'hd45f;
aud[9027]=16'hd46f;
aud[9028]=16'hd47f;
aud[9029]=16'hd48f;
aud[9030]=16'hd49e;
aud[9031]=16'hd4ae;
aud[9032]=16'hd4be;
aud[9033]=16'hd4ce;
aud[9034]=16'hd4de;
aud[9035]=16'hd4ed;
aud[9036]=16'hd4fd;
aud[9037]=16'hd50d;
aud[9038]=16'hd51d;
aud[9039]=16'hd52d;
aud[9040]=16'hd53d;
aud[9041]=16'hd54d;
aud[9042]=16'hd55d;
aud[9043]=16'hd56d;
aud[9044]=16'hd57d;
aud[9045]=16'hd58d;
aud[9046]=16'hd59d;
aud[9047]=16'hd5ad;
aud[9048]=16'hd5bd;
aud[9049]=16'hd5cd;
aud[9050]=16'hd5dd;
aud[9051]=16'hd5ee;
aud[9052]=16'hd5fe;
aud[9053]=16'hd60e;
aud[9054]=16'hd61e;
aud[9055]=16'hd62e;
aud[9056]=16'hd63f;
aud[9057]=16'hd64f;
aud[9058]=16'hd65f;
aud[9059]=16'hd66f;
aud[9060]=16'hd680;
aud[9061]=16'hd690;
aud[9062]=16'hd6a0;
aud[9063]=16'hd6b1;
aud[9064]=16'hd6c1;
aud[9065]=16'hd6d2;
aud[9066]=16'hd6e2;
aud[9067]=16'hd6f2;
aud[9068]=16'hd703;
aud[9069]=16'hd713;
aud[9070]=16'hd724;
aud[9071]=16'hd734;
aud[9072]=16'hd745;
aud[9073]=16'hd756;
aud[9074]=16'hd766;
aud[9075]=16'hd777;
aud[9076]=16'hd787;
aud[9077]=16'hd798;
aud[9078]=16'hd7a9;
aud[9079]=16'hd7b9;
aud[9080]=16'hd7ca;
aud[9081]=16'hd7db;
aud[9082]=16'hd7eb;
aud[9083]=16'hd7fc;
aud[9084]=16'hd80d;
aud[9085]=16'hd81e;
aud[9086]=16'hd82e;
aud[9087]=16'hd83f;
aud[9088]=16'hd850;
aud[9089]=16'hd861;
aud[9090]=16'hd872;
aud[9091]=16'hd882;
aud[9092]=16'hd893;
aud[9093]=16'hd8a4;
aud[9094]=16'hd8b5;
aud[9095]=16'hd8c6;
aud[9096]=16'hd8d7;
aud[9097]=16'hd8e8;
aud[9098]=16'hd8f9;
aud[9099]=16'hd90a;
aud[9100]=16'hd91b;
aud[9101]=16'hd92c;
aud[9102]=16'hd93d;
aud[9103]=16'hd94e;
aud[9104]=16'hd95f;
aud[9105]=16'hd970;
aud[9106]=16'hd982;
aud[9107]=16'hd993;
aud[9108]=16'hd9a4;
aud[9109]=16'hd9b5;
aud[9110]=16'hd9c6;
aud[9111]=16'hd9d7;
aud[9112]=16'hd9e9;
aud[9113]=16'hd9fa;
aud[9114]=16'hda0b;
aud[9115]=16'hda1c;
aud[9116]=16'hda2e;
aud[9117]=16'hda3f;
aud[9118]=16'hda50;
aud[9119]=16'hda62;
aud[9120]=16'hda73;
aud[9121]=16'hda84;
aud[9122]=16'hda96;
aud[9123]=16'hdaa7;
aud[9124]=16'hdab9;
aud[9125]=16'hdaca;
aud[9126]=16'hdadc;
aud[9127]=16'hdaed;
aud[9128]=16'hdaff;
aud[9129]=16'hdb10;
aud[9130]=16'hdb22;
aud[9131]=16'hdb33;
aud[9132]=16'hdb45;
aud[9133]=16'hdb56;
aud[9134]=16'hdb68;
aud[9135]=16'hdb79;
aud[9136]=16'hdb8b;
aud[9137]=16'hdb9d;
aud[9138]=16'hdbae;
aud[9139]=16'hdbc0;
aud[9140]=16'hdbd2;
aud[9141]=16'hdbe3;
aud[9142]=16'hdbf5;
aud[9143]=16'hdc07;
aud[9144]=16'hdc19;
aud[9145]=16'hdc2a;
aud[9146]=16'hdc3c;
aud[9147]=16'hdc4e;
aud[9148]=16'hdc60;
aud[9149]=16'hdc72;
aud[9150]=16'hdc83;
aud[9151]=16'hdc95;
aud[9152]=16'hdca7;
aud[9153]=16'hdcb9;
aud[9154]=16'hdccb;
aud[9155]=16'hdcdd;
aud[9156]=16'hdcef;
aud[9157]=16'hdd01;
aud[9158]=16'hdd13;
aud[9159]=16'hdd25;
aud[9160]=16'hdd37;
aud[9161]=16'hdd49;
aud[9162]=16'hdd5b;
aud[9163]=16'hdd6d;
aud[9164]=16'hdd7f;
aud[9165]=16'hdd91;
aud[9166]=16'hdda3;
aud[9167]=16'hddb5;
aud[9168]=16'hddc7;
aud[9169]=16'hddd9;
aud[9170]=16'hddeb;
aud[9171]=16'hddfe;
aud[9172]=16'hde10;
aud[9173]=16'hde22;
aud[9174]=16'hde34;
aud[9175]=16'hde46;
aud[9176]=16'hde59;
aud[9177]=16'hde6b;
aud[9178]=16'hde7d;
aud[9179]=16'hde8f;
aud[9180]=16'hdea2;
aud[9181]=16'hdeb4;
aud[9182]=16'hdec6;
aud[9183]=16'hded9;
aud[9184]=16'hdeeb;
aud[9185]=16'hdefd;
aud[9186]=16'hdf10;
aud[9187]=16'hdf22;
aud[9188]=16'hdf35;
aud[9189]=16'hdf47;
aud[9190]=16'hdf59;
aud[9191]=16'hdf6c;
aud[9192]=16'hdf7e;
aud[9193]=16'hdf91;
aud[9194]=16'hdfa3;
aud[9195]=16'hdfb6;
aud[9196]=16'hdfc8;
aud[9197]=16'hdfdb;
aud[9198]=16'hdfed;
aud[9199]=16'he000;
aud[9200]=16'he013;
aud[9201]=16'he025;
aud[9202]=16'he038;
aud[9203]=16'he04a;
aud[9204]=16'he05d;
aud[9205]=16'he070;
aud[9206]=16'he082;
aud[9207]=16'he095;
aud[9208]=16'he0a8;
aud[9209]=16'he0ba;
aud[9210]=16'he0cd;
aud[9211]=16'he0e0;
aud[9212]=16'he0f3;
aud[9213]=16'he105;
aud[9214]=16'he118;
aud[9215]=16'he12b;
aud[9216]=16'he13e;
aud[9217]=16'he151;
aud[9218]=16'he163;
aud[9219]=16'he176;
aud[9220]=16'he189;
aud[9221]=16'he19c;
aud[9222]=16'he1af;
aud[9223]=16'he1c2;
aud[9224]=16'he1d5;
aud[9225]=16'he1e8;
aud[9226]=16'he1fa;
aud[9227]=16'he20d;
aud[9228]=16'he220;
aud[9229]=16'he233;
aud[9230]=16'he246;
aud[9231]=16'he259;
aud[9232]=16'he26c;
aud[9233]=16'he27f;
aud[9234]=16'he292;
aud[9235]=16'he2a5;
aud[9236]=16'he2b9;
aud[9237]=16'he2cc;
aud[9238]=16'he2df;
aud[9239]=16'he2f2;
aud[9240]=16'he305;
aud[9241]=16'he318;
aud[9242]=16'he32b;
aud[9243]=16'he33e;
aud[9244]=16'he352;
aud[9245]=16'he365;
aud[9246]=16'he378;
aud[9247]=16'he38b;
aud[9248]=16'he39e;
aud[9249]=16'he3b2;
aud[9250]=16'he3c5;
aud[9251]=16'he3d8;
aud[9252]=16'he3eb;
aud[9253]=16'he3ff;
aud[9254]=16'he412;
aud[9255]=16'he425;
aud[9256]=16'he438;
aud[9257]=16'he44c;
aud[9258]=16'he45f;
aud[9259]=16'he473;
aud[9260]=16'he486;
aud[9261]=16'he499;
aud[9262]=16'he4ad;
aud[9263]=16'he4c0;
aud[9264]=16'he4d3;
aud[9265]=16'he4e7;
aud[9266]=16'he4fa;
aud[9267]=16'he50e;
aud[9268]=16'he521;
aud[9269]=16'he535;
aud[9270]=16'he548;
aud[9271]=16'he55c;
aud[9272]=16'he56f;
aud[9273]=16'he583;
aud[9274]=16'he596;
aud[9275]=16'he5aa;
aud[9276]=16'he5bd;
aud[9277]=16'he5d1;
aud[9278]=16'he5e4;
aud[9279]=16'he5f8;
aud[9280]=16'he60c;
aud[9281]=16'he61f;
aud[9282]=16'he633;
aud[9283]=16'he646;
aud[9284]=16'he65a;
aud[9285]=16'he66e;
aud[9286]=16'he681;
aud[9287]=16'he695;
aud[9288]=16'he6a9;
aud[9289]=16'he6bd;
aud[9290]=16'he6d0;
aud[9291]=16'he6e4;
aud[9292]=16'he6f8;
aud[9293]=16'he70b;
aud[9294]=16'he71f;
aud[9295]=16'he733;
aud[9296]=16'he747;
aud[9297]=16'he75b;
aud[9298]=16'he76e;
aud[9299]=16'he782;
aud[9300]=16'he796;
aud[9301]=16'he7aa;
aud[9302]=16'he7be;
aud[9303]=16'he7d1;
aud[9304]=16'he7e5;
aud[9305]=16'he7f9;
aud[9306]=16'he80d;
aud[9307]=16'he821;
aud[9308]=16'he835;
aud[9309]=16'he849;
aud[9310]=16'he85d;
aud[9311]=16'he871;
aud[9312]=16'he885;
aud[9313]=16'he899;
aud[9314]=16'he8ad;
aud[9315]=16'he8c0;
aud[9316]=16'he8d4;
aud[9317]=16'he8e8;
aud[9318]=16'he8fc;
aud[9319]=16'he910;
aud[9320]=16'he925;
aud[9321]=16'he939;
aud[9322]=16'he94d;
aud[9323]=16'he961;
aud[9324]=16'he975;
aud[9325]=16'he989;
aud[9326]=16'he99d;
aud[9327]=16'he9b1;
aud[9328]=16'he9c5;
aud[9329]=16'he9d9;
aud[9330]=16'he9ed;
aud[9331]=16'hea01;
aud[9332]=16'hea16;
aud[9333]=16'hea2a;
aud[9334]=16'hea3e;
aud[9335]=16'hea52;
aud[9336]=16'hea66;
aud[9337]=16'hea7a;
aud[9338]=16'hea8f;
aud[9339]=16'heaa3;
aud[9340]=16'heab7;
aud[9341]=16'heacb;
aud[9342]=16'heae0;
aud[9343]=16'heaf4;
aud[9344]=16'heb08;
aud[9345]=16'heb1c;
aud[9346]=16'heb31;
aud[9347]=16'heb45;
aud[9348]=16'heb59;
aud[9349]=16'heb6e;
aud[9350]=16'heb82;
aud[9351]=16'heb96;
aud[9352]=16'hebab;
aud[9353]=16'hebbf;
aud[9354]=16'hebd3;
aud[9355]=16'hebe8;
aud[9356]=16'hebfc;
aud[9357]=16'hec10;
aud[9358]=16'hec25;
aud[9359]=16'hec39;
aud[9360]=16'hec4d;
aud[9361]=16'hec62;
aud[9362]=16'hec76;
aud[9363]=16'hec8b;
aud[9364]=16'hec9f;
aud[9365]=16'hecb4;
aud[9366]=16'hecc8;
aud[9367]=16'hecdd;
aud[9368]=16'hecf1;
aud[9369]=16'hed05;
aud[9370]=16'hed1a;
aud[9371]=16'hed2e;
aud[9372]=16'hed43;
aud[9373]=16'hed57;
aud[9374]=16'hed6c;
aud[9375]=16'hed81;
aud[9376]=16'hed95;
aud[9377]=16'hedaa;
aud[9378]=16'hedbe;
aud[9379]=16'hedd3;
aud[9380]=16'hede7;
aud[9381]=16'hedfc;
aud[9382]=16'hee10;
aud[9383]=16'hee25;
aud[9384]=16'hee3a;
aud[9385]=16'hee4e;
aud[9386]=16'hee63;
aud[9387]=16'hee77;
aud[9388]=16'hee8c;
aud[9389]=16'heea1;
aud[9390]=16'heeb5;
aud[9391]=16'heeca;
aud[9392]=16'heedf;
aud[9393]=16'heef3;
aud[9394]=16'hef08;
aud[9395]=16'hef1d;
aud[9396]=16'hef31;
aud[9397]=16'hef46;
aud[9398]=16'hef5b;
aud[9399]=16'hef70;
aud[9400]=16'hef84;
aud[9401]=16'hef99;
aud[9402]=16'hefae;
aud[9403]=16'hefc2;
aud[9404]=16'hefd7;
aud[9405]=16'hefec;
aud[9406]=16'hf001;
aud[9407]=16'hf015;
aud[9408]=16'hf02a;
aud[9409]=16'hf03f;
aud[9410]=16'hf054;
aud[9411]=16'hf069;
aud[9412]=16'hf07d;
aud[9413]=16'hf092;
aud[9414]=16'hf0a7;
aud[9415]=16'hf0bc;
aud[9416]=16'hf0d1;
aud[9417]=16'hf0e6;
aud[9418]=16'hf0fa;
aud[9419]=16'hf10f;
aud[9420]=16'hf124;
aud[9421]=16'hf139;
aud[9422]=16'hf14e;
aud[9423]=16'hf163;
aud[9424]=16'hf178;
aud[9425]=16'hf18c;
aud[9426]=16'hf1a1;
aud[9427]=16'hf1b6;
aud[9428]=16'hf1cb;
aud[9429]=16'hf1e0;
aud[9430]=16'hf1f5;
aud[9431]=16'hf20a;
aud[9432]=16'hf21f;
aud[9433]=16'hf234;
aud[9434]=16'hf249;
aud[9435]=16'hf25e;
aud[9436]=16'hf273;
aud[9437]=16'hf288;
aud[9438]=16'hf29d;
aud[9439]=16'hf2b2;
aud[9440]=16'hf2c7;
aud[9441]=16'hf2dc;
aud[9442]=16'hf2f1;
aud[9443]=16'hf306;
aud[9444]=16'hf31b;
aud[9445]=16'hf330;
aud[9446]=16'hf345;
aud[9447]=16'hf35a;
aud[9448]=16'hf36f;
aud[9449]=16'hf384;
aud[9450]=16'hf399;
aud[9451]=16'hf3ae;
aud[9452]=16'hf3c3;
aud[9453]=16'hf3d8;
aud[9454]=16'hf3ed;
aud[9455]=16'hf402;
aud[9456]=16'hf417;
aud[9457]=16'hf42c;
aud[9458]=16'hf441;
aud[9459]=16'hf456;
aud[9460]=16'hf46b;
aud[9461]=16'hf480;
aud[9462]=16'hf496;
aud[9463]=16'hf4ab;
aud[9464]=16'hf4c0;
aud[9465]=16'hf4d5;
aud[9466]=16'hf4ea;
aud[9467]=16'hf4ff;
aud[9468]=16'hf514;
aud[9469]=16'hf529;
aud[9470]=16'hf53f;
aud[9471]=16'hf554;
aud[9472]=16'hf569;
aud[9473]=16'hf57e;
aud[9474]=16'hf593;
aud[9475]=16'hf5a8;
aud[9476]=16'hf5bd;
aud[9477]=16'hf5d3;
aud[9478]=16'hf5e8;
aud[9479]=16'hf5fd;
aud[9480]=16'hf612;
aud[9481]=16'hf627;
aud[9482]=16'hf63d;
aud[9483]=16'hf652;
aud[9484]=16'hf667;
aud[9485]=16'hf67c;
aud[9486]=16'hf691;
aud[9487]=16'hf6a7;
aud[9488]=16'hf6bc;
aud[9489]=16'hf6d1;
aud[9490]=16'hf6e6;
aud[9491]=16'hf6fb;
aud[9492]=16'hf711;
aud[9493]=16'hf726;
aud[9494]=16'hf73b;
aud[9495]=16'hf750;
aud[9496]=16'hf766;
aud[9497]=16'hf77b;
aud[9498]=16'hf790;
aud[9499]=16'hf7a5;
aud[9500]=16'hf7bb;
aud[9501]=16'hf7d0;
aud[9502]=16'hf7e5;
aud[9503]=16'hf7fb;
aud[9504]=16'hf810;
aud[9505]=16'hf825;
aud[9506]=16'hf83a;
aud[9507]=16'hf850;
aud[9508]=16'hf865;
aud[9509]=16'hf87a;
aud[9510]=16'hf890;
aud[9511]=16'hf8a5;
aud[9512]=16'hf8ba;
aud[9513]=16'hf8cf;
aud[9514]=16'hf8e5;
aud[9515]=16'hf8fa;
aud[9516]=16'hf90f;
aud[9517]=16'hf925;
aud[9518]=16'hf93a;
aud[9519]=16'hf94f;
aud[9520]=16'hf965;
aud[9521]=16'hf97a;
aud[9522]=16'hf98f;
aud[9523]=16'hf9a5;
aud[9524]=16'hf9ba;
aud[9525]=16'hf9cf;
aud[9526]=16'hf9e5;
aud[9527]=16'hf9fa;
aud[9528]=16'hfa0f;
aud[9529]=16'hfa25;
aud[9530]=16'hfa3a;
aud[9531]=16'hfa50;
aud[9532]=16'hfa65;
aud[9533]=16'hfa7a;
aud[9534]=16'hfa90;
aud[9535]=16'hfaa5;
aud[9536]=16'hfaba;
aud[9537]=16'hfad0;
aud[9538]=16'hfae5;
aud[9539]=16'hfafb;
aud[9540]=16'hfb10;
aud[9541]=16'hfb25;
aud[9542]=16'hfb3b;
aud[9543]=16'hfb50;
aud[9544]=16'hfb65;
aud[9545]=16'hfb7b;
aud[9546]=16'hfb90;
aud[9547]=16'hfba6;
aud[9548]=16'hfbbb;
aud[9549]=16'hfbd0;
aud[9550]=16'hfbe6;
aud[9551]=16'hfbfb;
aud[9552]=16'hfc11;
aud[9553]=16'hfc26;
aud[9554]=16'hfc3b;
aud[9555]=16'hfc51;
aud[9556]=16'hfc66;
aud[9557]=16'hfc7c;
aud[9558]=16'hfc91;
aud[9559]=16'hfca7;
aud[9560]=16'hfcbc;
aud[9561]=16'hfcd1;
aud[9562]=16'hfce7;
aud[9563]=16'hfcfc;
aud[9564]=16'hfd12;
aud[9565]=16'hfd27;
aud[9566]=16'hfd3c;
aud[9567]=16'hfd52;
aud[9568]=16'hfd67;
aud[9569]=16'hfd7d;
aud[9570]=16'hfd92;
aud[9571]=16'hfda8;
aud[9572]=16'hfdbd;
aud[9573]=16'hfdd2;
aud[9574]=16'hfde8;
aud[9575]=16'hfdfd;
aud[9576]=16'hfe13;
aud[9577]=16'hfe28;
aud[9578]=16'hfe3e;
aud[9579]=16'hfe53;
aud[9580]=16'hfe69;
aud[9581]=16'hfe7e;
aud[9582]=16'hfe93;
aud[9583]=16'hfea9;
aud[9584]=16'hfebe;
aud[9585]=16'hfed4;
aud[9586]=16'hfee9;
aud[9587]=16'hfeff;
aud[9588]=16'hff14;
aud[9589]=16'hff2a;
aud[9590]=16'hff3f;
aud[9591]=16'hff54;
aud[9592]=16'hff6a;
aud[9593]=16'hff7f;
aud[9594]=16'hff95;
aud[9595]=16'hffaa;
aud[9596]=16'hffc0;
aud[9597]=16'hffd5;
aud[9598]=16'hffeb;
aud[9599]=16'h0;
aud[9600]=16'h15;
aud[9601]=16'h2b;
aud[9602]=16'h40;
aud[9603]=16'h56;
aud[9604]=16'h6b;
aud[9605]=16'h81;
aud[9606]=16'h96;
aud[9607]=16'hac;
aud[9608]=16'hc1;
aud[9609]=16'hd6;
aud[9610]=16'hec;
aud[9611]=16'h101;
aud[9612]=16'h117;
aud[9613]=16'h12c;
aud[9614]=16'h142;
aud[9615]=16'h157;
aud[9616]=16'h16d;
aud[9617]=16'h182;
aud[9618]=16'h197;
aud[9619]=16'h1ad;
aud[9620]=16'h1c2;
aud[9621]=16'h1d8;
aud[9622]=16'h1ed;
aud[9623]=16'h203;
aud[9624]=16'h218;
aud[9625]=16'h22e;
aud[9626]=16'h243;
aud[9627]=16'h258;
aud[9628]=16'h26e;
aud[9629]=16'h283;
aud[9630]=16'h299;
aud[9631]=16'h2ae;
aud[9632]=16'h2c4;
aud[9633]=16'h2d9;
aud[9634]=16'h2ee;
aud[9635]=16'h304;
aud[9636]=16'h319;
aud[9637]=16'h32f;
aud[9638]=16'h344;
aud[9639]=16'h359;
aud[9640]=16'h36f;
aud[9641]=16'h384;
aud[9642]=16'h39a;
aud[9643]=16'h3af;
aud[9644]=16'h3c5;
aud[9645]=16'h3da;
aud[9646]=16'h3ef;
aud[9647]=16'h405;
aud[9648]=16'h41a;
aud[9649]=16'h430;
aud[9650]=16'h445;
aud[9651]=16'h45a;
aud[9652]=16'h470;
aud[9653]=16'h485;
aud[9654]=16'h49b;
aud[9655]=16'h4b0;
aud[9656]=16'h4c5;
aud[9657]=16'h4db;
aud[9658]=16'h4f0;
aud[9659]=16'h505;
aud[9660]=16'h51b;
aud[9661]=16'h530;
aud[9662]=16'h546;
aud[9663]=16'h55b;
aud[9664]=16'h570;
aud[9665]=16'h586;
aud[9666]=16'h59b;
aud[9667]=16'h5b0;
aud[9668]=16'h5c6;
aud[9669]=16'h5db;
aud[9670]=16'h5f1;
aud[9671]=16'h606;
aud[9672]=16'h61b;
aud[9673]=16'h631;
aud[9674]=16'h646;
aud[9675]=16'h65b;
aud[9676]=16'h671;
aud[9677]=16'h686;
aud[9678]=16'h69b;
aud[9679]=16'h6b1;
aud[9680]=16'h6c6;
aud[9681]=16'h6db;
aud[9682]=16'h6f1;
aud[9683]=16'h706;
aud[9684]=16'h71b;
aud[9685]=16'h731;
aud[9686]=16'h746;
aud[9687]=16'h75b;
aud[9688]=16'h770;
aud[9689]=16'h786;
aud[9690]=16'h79b;
aud[9691]=16'h7b0;
aud[9692]=16'h7c6;
aud[9693]=16'h7db;
aud[9694]=16'h7f0;
aud[9695]=16'h805;
aud[9696]=16'h81b;
aud[9697]=16'h830;
aud[9698]=16'h845;
aud[9699]=16'h85b;
aud[9700]=16'h870;
aud[9701]=16'h885;
aud[9702]=16'h89a;
aud[9703]=16'h8b0;
aud[9704]=16'h8c5;
aud[9705]=16'h8da;
aud[9706]=16'h8ef;
aud[9707]=16'h905;
aud[9708]=16'h91a;
aud[9709]=16'h92f;
aud[9710]=16'h944;
aud[9711]=16'h959;
aud[9712]=16'h96f;
aud[9713]=16'h984;
aud[9714]=16'h999;
aud[9715]=16'h9ae;
aud[9716]=16'h9c3;
aud[9717]=16'h9d9;
aud[9718]=16'h9ee;
aud[9719]=16'ha03;
aud[9720]=16'ha18;
aud[9721]=16'ha2d;
aud[9722]=16'ha43;
aud[9723]=16'ha58;
aud[9724]=16'ha6d;
aud[9725]=16'ha82;
aud[9726]=16'ha97;
aud[9727]=16'haac;
aud[9728]=16'hac1;
aud[9729]=16'had7;
aud[9730]=16'haec;
aud[9731]=16'hb01;
aud[9732]=16'hb16;
aud[9733]=16'hb2b;
aud[9734]=16'hb40;
aud[9735]=16'hb55;
aud[9736]=16'hb6a;
aud[9737]=16'hb80;
aud[9738]=16'hb95;
aud[9739]=16'hbaa;
aud[9740]=16'hbbf;
aud[9741]=16'hbd4;
aud[9742]=16'hbe9;
aud[9743]=16'hbfe;
aud[9744]=16'hc13;
aud[9745]=16'hc28;
aud[9746]=16'hc3d;
aud[9747]=16'hc52;
aud[9748]=16'hc67;
aud[9749]=16'hc7c;
aud[9750]=16'hc91;
aud[9751]=16'hca6;
aud[9752]=16'hcbb;
aud[9753]=16'hcd0;
aud[9754]=16'hce5;
aud[9755]=16'hcfa;
aud[9756]=16'hd0f;
aud[9757]=16'hd24;
aud[9758]=16'hd39;
aud[9759]=16'hd4e;
aud[9760]=16'hd63;
aud[9761]=16'hd78;
aud[9762]=16'hd8d;
aud[9763]=16'hda2;
aud[9764]=16'hdb7;
aud[9765]=16'hdcc;
aud[9766]=16'hde1;
aud[9767]=16'hdf6;
aud[9768]=16'he0b;
aud[9769]=16'he20;
aud[9770]=16'he35;
aud[9771]=16'he4a;
aud[9772]=16'he5f;
aud[9773]=16'he74;
aud[9774]=16'he88;
aud[9775]=16'he9d;
aud[9776]=16'heb2;
aud[9777]=16'hec7;
aud[9778]=16'hedc;
aud[9779]=16'hef1;
aud[9780]=16'hf06;
aud[9781]=16'hf1a;
aud[9782]=16'hf2f;
aud[9783]=16'hf44;
aud[9784]=16'hf59;
aud[9785]=16'hf6e;
aud[9786]=16'hf83;
aud[9787]=16'hf97;
aud[9788]=16'hfac;
aud[9789]=16'hfc1;
aud[9790]=16'hfd6;
aud[9791]=16'hfeb;
aud[9792]=16'hfff;
aud[9793]=16'h1014;
aud[9794]=16'h1029;
aud[9795]=16'h103e;
aud[9796]=16'h1052;
aud[9797]=16'h1067;
aud[9798]=16'h107c;
aud[9799]=16'h1090;
aud[9800]=16'h10a5;
aud[9801]=16'h10ba;
aud[9802]=16'h10cf;
aud[9803]=16'h10e3;
aud[9804]=16'h10f8;
aud[9805]=16'h110d;
aud[9806]=16'h1121;
aud[9807]=16'h1136;
aud[9808]=16'h114b;
aud[9809]=16'h115f;
aud[9810]=16'h1174;
aud[9811]=16'h1189;
aud[9812]=16'h119d;
aud[9813]=16'h11b2;
aud[9814]=16'h11c6;
aud[9815]=16'h11db;
aud[9816]=16'h11f0;
aud[9817]=16'h1204;
aud[9818]=16'h1219;
aud[9819]=16'h122d;
aud[9820]=16'h1242;
aud[9821]=16'h1256;
aud[9822]=16'h126b;
aud[9823]=16'h127f;
aud[9824]=16'h1294;
aud[9825]=16'h12a9;
aud[9826]=16'h12bd;
aud[9827]=16'h12d2;
aud[9828]=16'h12e6;
aud[9829]=16'h12fb;
aud[9830]=16'h130f;
aud[9831]=16'h1323;
aud[9832]=16'h1338;
aud[9833]=16'h134c;
aud[9834]=16'h1361;
aud[9835]=16'h1375;
aud[9836]=16'h138a;
aud[9837]=16'h139e;
aud[9838]=16'h13b3;
aud[9839]=16'h13c7;
aud[9840]=16'h13db;
aud[9841]=16'h13f0;
aud[9842]=16'h1404;
aud[9843]=16'h1418;
aud[9844]=16'h142d;
aud[9845]=16'h1441;
aud[9846]=16'h1455;
aud[9847]=16'h146a;
aud[9848]=16'h147e;
aud[9849]=16'h1492;
aud[9850]=16'h14a7;
aud[9851]=16'h14bb;
aud[9852]=16'h14cf;
aud[9853]=16'h14e4;
aud[9854]=16'h14f8;
aud[9855]=16'h150c;
aud[9856]=16'h1520;
aud[9857]=16'h1535;
aud[9858]=16'h1549;
aud[9859]=16'h155d;
aud[9860]=16'h1571;
aud[9861]=16'h1586;
aud[9862]=16'h159a;
aud[9863]=16'h15ae;
aud[9864]=16'h15c2;
aud[9865]=16'h15d6;
aud[9866]=16'h15ea;
aud[9867]=16'h15ff;
aud[9868]=16'h1613;
aud[9869]=16'h1627;
aud[9870]=16'h163b;
aud[9871]=16'h164f;
aud[9872]=16'h1663;
aud[9873]=16'h1677;
aud[9874]=16'h168b;
aud[9875]=16'h169f;
aud[9876]=16'h16b3;
aud[9877]=16'h16c7;
aud[9878]=16'h16db;
aud[9879]=16'h16f0;
aud[9880]=16'h1704;
aud[9881]=16'h1718;
aud[9882]=16'h172c;
aud[9883]=16'h1740;
aud[9884]=16'h1753;
aud[9885]=16'h1767;
aud[9886]=16'h177b;
aud[9887]=16'h178f;
aud[9888]=16'h17a3;
aud[9889]=16'h17b7;
aud[9890]=16'h17cb;
aud[9891]=16'h17df;
aud[9892]=16'h17f3;
aud[9893]=16'h1807;
aud[9894]=16'h181b;
aud[9895]=16'h182f;
aud[9896]=16'h1842;
aud[9897]=16'h1856;
aud[9898]=16'h186a;
aud[9899]=16'h187e;
aud[9900]=16'h1892;
aud[9901]=16'h18a5;
aud[9902]=16'h18b9;
aud[9903]=16'h18cd;
aud[9904]=16'h18e1;
aud[9905]=16'h18f5;
aud[9906]=16'h1908;
aud[9907]=16'h191c;
aud[9908]=16'h1930;
aud[9909]=16'h1943;
aud[9910]=16'h1957;
aud[9911]=16'h196b;
aud[9912]=16'h197f;
aud[9913]=16'h1992;
aud[9914]=16'h19a6;
aud[9915]=16'h19ba;
aud[9916]=16'h19cd;
aud[9917]=16'h19e1;
aud[9918]=16'h19f4;
aud[9919]=16'h1a08;
aud[9920]=16'h1a1c;
aud[9921]=16'h1a2f;
aud[9922]=16'h1a43;
aud[9923]=16'h1a56;
aud[9924]=16'h1a6a;
aud[9925]=16'h1a7d;
aud[9926]=16'h1a91;
aud[9927]=16'h1aa4;
aud[9928]=16'h1ab8;
aud[9929]=16'h1acb;
aud[9930]=16'h1adf;
aud[9931]=16'h1af2;
aud[9932]=16'h1b06;
aud[9933]=16'h1b19;
aud[9934]=16'h1b2d;
aud[9935]=16'h1b40;
aud[9936]=16'h1b53;
aud[9937]=16'h1b67;
aud[9938]=16'h1b7a;
aud[9939]=16'h1b8d;
aud[9940]=16'h1ba1;
aud[9941]=16'h1bb4;
aud[9942]=16'h1bc8;
aud[9943]=16'h1bdb;
aud[9944]=16'h1bee;
aud[9945]=16'h1c01;
aud[9946]=16'h1c15;
aud[9947]=16'h1c28;
aud[9948]=16'h1c3b;
aud[9949]=16'h1c4e;
aud[9950]=16'h1c62;
aud[9951]=16'h1c75;
aud[9952]=16'h1c88;
aud[9953]=16'h1c9b;
aud[9954]=16'h1cae;
aud[9955]=16'h1cc2;
aud[9956]=16'h1cd5;
aud[9957]=16'h1ce8;
aud[9958]=16'h1cfb;
aud[9959]=16'h1d0e;
aud[9960]=16'h1d21;
aud[9961]=16'h1d34;
aud[9962]=16'h1d47;
aud[9963]=16'h1d5b;
aud[9964]=16'h1d6e;
aud[9965]=16'h1d81;
aud[9966]=16'h1d94;
aud[9967]=16'h1da7;
aud[9968]=16'h1dba;
aud[9969]=16'h1dcd;
aud[9970]=16'h1de0;
aud[9971]=16'h1df3;
aud[9972]=16'h1e06;
aud[9973]=16'h1e18;
aud[9974]=16'h1e2b;
aud[9975]=16'h1e3e;
aud[9976]=16'h1e51;
aud[9977]=16'h1e64;
aud[9978]=16'h1e77;
aud[9979]=16'h1e8a;
aud[9980]=16'h1e9d;
aud[9981]=16'h1eaf;
aud[9982]=16'h1ec2;
aud[9983]=16'h1ed5;
aud[9984]=16'h1ee8;
aud[9985]=16'h1efb;
aud[9986]=16'h1f0d;
aud[9987]=16'h1f20;
aud[9988]=16'h1f33;
aud[9989]=16'h1f46;
aud[9990]=16'h1f58;
aud[9991]=16'h1f6b;
aud[9992]=16'h1f7e;
aud[9993]=16'h1f90;
aud[9994]=16'h1fa3;
aud[9995]=16'h1fb6;
aud[9996]=16'h1fc8;
aud[9997]=16'h1fdb;
aud[9998]=16'h1fed;
aud[9999]=16'h2000;
aud[10000]=16'h2013;
aud[10001]=16'h2025;
aud[10002]=16'h2038;
aud[10003]=16'h204a;
aud[10004]=16'h205d;
aud[10005]=16'h206f;
aud[10006]=16'h2082;
aud[10007]=16'h2094;
aud[10008]=16'h20a7;
aud[10009]=16'h20b9;
aud[10010]=16'h20cb;
aud[10011]=16'h20de;
aud[10012]=16'h20f0;
aud[10013]=16'h2103;
aud[10014]=16'h2115;
aud[10015]=16'h2127;
aud[10016]=16'h213a;
aud[10017]=16'h214c;
aud[10018]=16'h215e;
aud[10019]=16'h2171;
aud[10020]=16'h2183;
aud[10021]=16'h2195;
aud[10022]=16'h21a7;
aud[10023]=16'h21ba;
aud[10024]=16'h21cc;
aud[10025]=16'h21de;
aud[10026]=16'h21f0;
aud[10027]=16'h2202;
aud[10028]=16'h2215;
aud[10029]=16'h2227;
aud[10030]=16'h2239;
aud[10031]=16'h224b;
aud[10032]=16'h225d;
aud[10033]=16'h226f;
aud[10034]=16'h2281;
aud[10035]=16'h2293;
aud[10036]=16'h22a5;
aud[10037]=16'h22b7;
aud[10038]=16'h22c9;
aud[10039]=16'h22db;
aud[10040]=16'h22ed;
aud[10041]=16'h22ff;
aud[10042]=16'h2311;
aud[10043]=16'h2323;
aud[10044]=16'h2335;
aud[10045]=16'h2347;
aud[10046]=16'h2359;
aud[10047]=16'h236b;
aud[10048]=16'h237d;
aud[10049]=16'h238e;
aud[10050]=16'h23a0;
aud[10051]=16'h23b2;
aud[10052]=16'h23c4;
aud[10053]=16'h23d6;
aud[10054]=16'h23e7;
aud[10055]=16'h23f9;
aud[10056]=16'h240b;
aud[10057]=16'h241d;
aud[10058]=16'h242e;
aud[10059]=16'h2440;
aud[10060]=16'h2452;
aud[10061]=16'h2463;
aud[10062]=16'h2475;
aud[10063]=16'h2487;
aud[10064]=16'h2498;
aud[10065]=16'h24aa;
aud[10066]=16'h24bb;
aud[10067]=16'h24cd;
aud[10068]=16'h24de;
aud[10069]=16'h24f0;
aud[10070]=16'h2501;
aud[10071]=16'h2513;
aud[10072]=16'h2524;
aud[10073]=16'h2536;
aud[10074]=16'h2547;
aud[10075]=16'h2559;
aud[10076]=16'h256a;
aud[10077]=16'h257c;
aud[10078]=16'h258d;
aud[10079]=16'h259e;
aud[10080]=16'h25b0;
aud[10081]=16'h25c1;
aud[10082]=16'h25d2;
aud[10083]=16'h25e4;
aud[10084]=16'h25f5;
aud[10085]=16'h2606;
aud[10086]=16'h2617;
aud[10087]=16'h2629;
aud[10088]=16'h263a;
aud[10089]=16'h264b;
aud[10090]=16'h265c;
aud[10091]=16'h266d;
aud[10092]=16'h267e;
aud[10093]=16'h2690;
aud[10094]=16'h26a1;
aud[10095]=16'h26b2;
aud[10096]=16'h26c3;
aud[10097]=16'h26d4;
aud[10098]=16'h26e5;
aud[10099]=16'h26f6;
aud[10100]=16'h2707;
aud[10101]=16'h2718;
aud[10102]=16'h2729;
aud[10103]=16'h273a;
aud[10104]=16'h274b;
aud[10105]=16'h275c;
aud[10106]=16'h276d;
aud[10107]=16'h277e;
aud[10108]=16'h278e;
aud[10109]=16'h279f;
aud[10110]=16'h27b0;
aud[10111]=16'h27c1;
aud[10112]=16'h27d2;
aud[10113]=16'h27e2;
aud[10114]=16'h27f3;
aud[10115]=16'h2804;
aud[10116]=16'h2815;
aud[10117]=16'h2825;
aud[10118]=16'h2836;
aud[10119]=16'h2847;
aud[10120]=16'h2857;
aud[10121]=16'h2868;
aud[10122]=16'h2879;
aud[10123]=16'h2889;
aud[10124]=16'h289a;
aud[10125]=16'h28aa;
aud[10126]=16'h28bb;
aud[10127]=16'h28cc;
aud[10128]=16'h28dc;
aud[10129]=16'h28ed;
aud[10130]=16'h28fd;
aud[10131]=16'h290e;
aud[10132]=16'h291e;
aud[10133]=16'h292e;
aud[10134]=16'h293f;
aud[10135]=16'h294f;
aud[10136]=16'h2960;
aud[10137]=16'h2970;
aud[10138]=16'h2980;
aud[10139]=16'h2991;
aud[10140]=16'h29a1;
aud[10141]=16'h29b1;
aud[10142]=16'h29c1;
aud[10143]=16'h29d2;
aud[10144]=16'h29e2;
aud[10145]=16'h29f2;
aud[10146]=16'h2a02;
aud[10147]=16'h2a12;
aud[10148]=16'h2a23;
aud[10149]=16'h2a33;
aud[10150]=16'h2a43;
aud[10151]=16'h2a53;
aud[10152]=16'h2a63;
aud[10153]=16'h2a73;
aud[10154]=16'h2a83;
aud[10155]=16'h2a93;
aud[10156]=16'h2aa3;
aud[10157]=16'h2ab3;
aud[10158]=16'h2ac3;
aud[10159]=16'h2ad3;
aud[10160]=16'h2ae3;
aud[10161]=16'h2af3;
aud[10162]=16'h2b03;
aud[10163]=16'h2b13;
aud[10164]=16'h2b22;
aud[10165]=16'h2b32;
aud[10166]=16'h2b42;
aud[10167]=16'h2b52;
aud[10168]=16'h2b62;
aud[10169]=16'h2b71;
aud[10170]=16'h2b81;
aud[10171]=16'h2b91;
aud[10172]=16'h2ba1;
aud[10173]=16'h2bb0;
aud[10174]=16'h2bc0;
aud[10175]=16'h2bd0;
aud[10176]=16'h2bdf;
aud[10177]=16'h2bef;
aud[10178]=16'h2bfe;
aud[10179]=16'h2c0e;
aud[10180]=16'h2c1e;
aud[10181]=16'h2c2d;
aud[10182]=16'h2c3d;
aud[10183]=16'h2c4c;
aud[10184]=16'h2c5c;
aud[10185]=16'h2c6b;
aud[10186]=16'h2c7a;
aud[10187]=16'h2c8a;
aud[10188]=16'h2c99;
aud[10189]=16'h2ca9;
aud[10190]=16'h2cb8;
aud[10191]=16'h2cc7;
aud[10192]=16'h2cd7;
aud[10193]=16'h2ce6;
aud[10194]=16'h2cf5;
aud[10195]=16'h2d04;
aud[10196]=16'h2d14;
aud[10197]=16'h2d23;
aud[10198]=16'h2d32;
aud[10199]=16'h2d41;
aud[10200]=16'h2d50;
aud[10201]=16'h2d60;
aud[10202]=16'h2d6f;
aud[10203]=16'h2d7e;
aud[10204]=16'h2d8d;
aud[10205]=16'h2d9c;
aud[10206]=16'h2dab;
aud[10207]=16'h2dba;
aud[10208]=16'h2dc9;
aud[10209]=16'h2dd8;
aud[10210]=16'h2de7;
aud[10211]=16'h2df6;
aud[10212]=16'h2e05;
aud[10213]=16'h2e14;
aud[10214]=16'h2e22;
aud[10215]=16'h2e31;
aud[10216]=16'h2e40;
aud[10217]=16'h2e4f;
aud[10218]=16'h2e5e;
aud[10219]=16'h2e6d;
aud[10220]=16'h2e7b;
aud[10221]=16'h2e8a;
aud[10222]=16'h2e99;
aud[10223]=16'h2ea7;
aud[10224]=16'h2eb6;
aud[10225]=16'h2ec5;
aud[10226]=16'h2ed3;
aud[10227]=16'h2ee2;
aud[10228]=16'h2ef1;
aud[10229]=16'h2eff;
aud[10230]=16'h2f0e;
aud[10231]=16'h2f1c;
aud[10232]=16'h2f2b;
aud[10233]=16'h2f39;
aud[10234]=16'h2f48;
aud[10235]=16'h2f56;
aud[10236]=16'h2f65;
aud[10237]=16'h2f73;
aud[10238]=16'h2f81;
aud[10239]=16'h2f90;
aud[10240]=16'h2f9e;
aud[10241]=16'h2fac;
aud[10242]=16'h2fbb;
aud[10243]=16'h2fc9;
aud[10244]=16'h2fd7;
aud[10245]=16'h2fe5;
aud[10246]=16'h2ff4;
aud[10247]=16'h3002;
aud[10248]=16'h3010;
aud[10249]=16'h301e;
aud[10250]=16'h302c;
aud[10251]=16'h303a;
aud[10252]=16'h3048;
aud[10253]=16'h3057;
aud[10254]=16'h3065;
aud[10255]=16'h3073;
aud[10256]=16'h3081;
aud[10257]=16'h308f;
aud[10258]=16'h309d;
aud[10259]=16'h30aa;
aud[10260]=16'h30b8;
aud[10261]=16'h30c6;
aud[10262]=16'h30d4;
aud[10263]=16'h30e2;
aud[10264]=16'h30f0;
aud[10265]=16'h30fe;
aud[10266]=16'h310b;
aud[10267]=16'h3119;
aud[10268]=16'h3127;
aud[10269]=16'h3135;
aud[10270]=16'h3142;
aud[10271]=16'h3150;
aud[10272]=16'h315e;
aud[10273]=16'h316b;
aud[10274]=16'h3179;
aud[10275]=16'h3187;
aud[10276]=16'h3194;
aud[10277]=16'h31a2;
aud[10278]=16'h31af;
aud[10279]=16'h31bd;
aud[10280]=16'h31ca;
aud[10281]=16'h31d8;
aud[10282]=16'h31e5;
aud[10283]=16'h31f3;
aud[10284]=16'h3200;
aud[10285]=16'h320d;
aud[10286]=16'h321b;
aud[10287]=16'h3228;
aud[10288]=16'h3235;
aud[10289]=16'h3243;
aud[10290]=16'h3250;
aud[10291]=16'h325d;
aud[10292]=16'h326a;
aud[10293]=16'h3278;
aud[10294]=16'h3285;
aud[10295]=16'h3292;
aud[10296]=16'h329f;
aud[10297]=16'h32ac;
aud[10298]=16'h32b9;
aud[10299]=16'h32c6;
aud[10300]=16'h32d3;
aud[10301]=16'h32e0;
aud[10302]=16'h32ed;
aud[10303]=16'h32fa;
aud[10304]=16'h3307;
aud[10305]=16'h3314;
aud[10306]=16'h3321;
aud[10307]=16'h332e;
aud[10308]=16'h333b;
aud[10309]=16'h3348;
aud[10310]=16'h3355;
aud[10311]=16'h3361;
aud[10312]=16'h336e;
aud[10313]=16'h337b;
aud[10314]=16'h3388;
aud[10315]=16'h3394;
aud[10316]=16'h33a1;
aud[10317]=16'h33ae;
aud[10318]=16'h33ba;
aud[10319]=16'h33c7;
aud[10320]=16'h33d4;
aud[10321]=16'h33e0;
aud[10322]=16'h33ed;
aud[10323]=16'h33f9;
aud[10324]=16'h3406;
aud[10325]=16'h3412;
aud[10326]=16'h341f;
aud[10327]=16'h342b;
aud[10328]=16'h3437;
aud[10329]=16'h3444;
aud[10330]=16'h3450;
aud[10331]=16'h345d;
aud[10332]=16'h3469;
aud[10333]=16'h3475;
aud[10334]=16'h3481;
aud[10335]=16'h348e;
aud[10336]=16'h349a;
aud[10337]=16'h34a6;
aud[10338]=16'h34b2;
aud[10339]=16'h34be;
aud[10340]=16'h34cb;
aud[10341]=16'h34d7;
aud[10342]=16'h34e3;
aud[10343]=16'h34ef;
aud[10344]=16'h34fb;
aud[10345]=16'h3507;
aud[10346]=16'h3513;
aud[10347]=16'h351f;
aud[10348]=16'h352b;
aud[10349]=16'h3537;
aud[10350]=16'h3543;
aud[10351]=16'h354f;
aud[10352]=16'h355a;
aud[10353]=16'h3566;
aud[10354]=16'h3572;
aud[10355]=16'h357e;
aud[10356]=16'h358a;
aud[10357]=16'h3595;
aud[10358]=16'h35a1;
aud[10359]=16'h35ad;
aud[10360]=16'h35b8;
aud[10361]=16'h35c4;
aud[10362]=16'h35d0;
aud[10363]=16'h35db;
aud[10364]=16'h35e7;
aud[10365]=16'h35f2;
aud[10366]=16'h35fe;
aud[10367]=16'h3609;
aud[10368]=16'h3615;
aud[10369]=16'h3620;
aud[10370]=16'h362c;
aud[10371]=16'h3637;
aud[10372]=16'h3643;
aud[10373]=16'h364e;
aud[10374]=16'h3659;
aud[10375]=16'h3665;
aud[10376]=16'h3670;
aud[10377]=16'h367b;
aud[10378]=16'h3686;
aud[10379]=16'h3692;
aud[10380]=16'h369d;
aud[10381]=16'h36a8;
aud[10382]=16'h36b3;
aud[10383]=16'h36be;
aud[10384]=16'h36c9;
aud[10385]=16'h36d4;
aud[10386]=16'h36e0;
aud[10387]=16'h36eb;
aud[10388]=16'h36f6;
aud[10389]=16'h3701;
aud[10390]=16'h370b;
aud[10391]=16'h3716;
aud[10392]=16'h3721;
aud[10393]=16'h372c;
aud[10394]=16'h3737;
aud[10395]=16'h3742;
aud[10396]=16'h374d;
aud[10397]=16'h3757;
aud[10398]=16'h3762;
aud[10399]=16'h376d;
aud[10400]=16'h3778;
aud[10401]=16'h3782;
aud[10402]=16'h378d;
aud[10403]=16'h3798;
aud[10404]=16'h37a2;
aud[10405]=16'h37ad;
aud[10406]=16'h37b7;
aud[10407]=16'h37c2;
aud[10408]=16'h37cc;
aud[10409]=16'h37d7;
aud[10410]=16'h37e1;
aud[10411]=16'h37ec;
aud[10412]=16'h37f6;
aud[10413]=16'h3801;
aud[10414]=16'h380b;
aud[10415]=16'h3815;
aud[10416]=16'h3820;
aud[10417]=16'h382a;
aud[10418]=16'h3834;
aud[10419]=16'h383f;
aud[10420]=16'h3849;
aud[10421]=16'h3853;
aud[10422]=16'h385d;
aud[10423]=16'h3867;
aud[10424]=16'h3871;
aud[10425]=16'h387b;
aud[10426]=16'h3886;
aud[10427]=16'h3890;
aud[10428]=16'h389a;
aud[10429]=16'h38a4;
aud[10430]=16'h38ae;
aud[10431]=16'h38b8;
aud[10432]=16'h38c1;
aud[10433]=16'h38cb;
aud[10434]=16'h38d5;
aud[10435]=16'h38df;
aud[10436]=16'h38e9;
aud[10437]=16'h38f3;
aud[10438]=16'h38fd;
aud[10439]=16'h3906;
aud[10440]=16'h3910;
aud[10441]=16'h391a;
aud[10442]=16'h3923;
aud[10443]=16'h392d;
aud[10444]=16'h3937;
aud[10445]=16'h3940;
aud[10446]=16'h394a;
aud[10447]=16'h3953;
aud[10448]=16'h395d;
aud[10449]=16'h3966;
aud[10450]=16'h3970;
aud[10451]=16'h3979;
aud[10452]=16'h3983;
aud[10453]=16'h398c;
aud[10454]=16'h3995;
aud[10455]=16'h399f;
aud[10456]=16'h39a8;
aud[10457]=16'h39b1;
aud[10458]=16'h39bb;
aud[10459]=16'h39c4;
aud[10460]=16'h39cd;
aud[10461]=16'h39d6;
aud[10462]=16'h39e0;
aud[10463]=16'h39e9;
aud[10464]=16'h39f2;
aud[10465]=16'h39fb;
aud[10466]=16'h3a04;
aud[10467]=16'h3a0d;
aud[10468]=16'h3a16;
aud[10469]=16'h3a1f;
aud[10470]=16'h3a28;
aud[10471]=16'h3a31;
aud[10472]=16'h3a3a;
aud[10473]=16'h3a43;
aud[10474]=16'h3a4c;
aud[10475]=16'h3a54;
aud[10476]=16'h3a5d;
aud[10477]=16'h3a66;
aud[10478]=16'h3a6f;
aud[10479]=16'h3a78;
aud[10480]=16'h3a80;
aud[10481]=16'h3a89;
aud[10482]=16'h3a92;
aud[10483]=16'h3a9a;
aud[10484]=16'h3aa3;
aud[10485]=16'h3aab;
aud[10486]=16'h3ab4;
aud[10487]=16'h3abc;
aud[10488]=16'h3ac5;
aud[10489]=16'h3acd;
aud[10490]=16'h3ad6;
aud[10491]=16'h3ade;
aud[10492]=16'h3ae7;
aud[10493]=16'h3aef;
aud[10494]=16'h3af7;
aud[10495]=16'h3b00;
aud[10496]=16'h3b08;
aud[10497]=16'h3b10;
aud[10498]=16'h3b19;
aud[10499]=16'h3b21;
aud[10500]=16'h3b29;
aud[10501]=16'h3b31;
aud[10502]=16'h3b39;
aud[10503]=16'h3b41;
aud[10504]=16'h3b4a;
aud[10505]=16'h3b52;
aud[10506]=16'h3b5a;
aud[10507]=16'h3b62;
aud[10508]=16'h3b6a;
aud[10509]=16'h3b72;
aud[10510]=16'h3b7a;
aud[10511]=16'h3b81;
aud[10512]=16'h3b89;
aud[10513]=16'h3b91;
aud[10514]=16'h3b99;
aud[10515]=16'h3ba1;
aud[10516]=16'h3ba9;
aud[10517]=16'h3bb0;
aud[10518]=16'h3bb8;
aud[10519]=16'h3bc0;
aud[10520]=16'h3bc7;
aud[10521]=16'h3bcf;
aud[10522]=16'h3bd7;
aud[10523]=16'h3bde;
aud[10524]=16'h3be6;
aud[10525]=16'h3bed;
aud[10526]=16'h3bf5;
aud[10527]=16'h3bfc;
aud[10528]=16'h3c04;
aud[10529]=16'h3c0b;
aud[10530]=16'h3c13;
aud[10531]=16'h3c1a;
aud[10532]=16'h3c21;
aud[10533]=16'h3c29;
aud[10534]=16'h3c30;
aud[10535]=16'h3c37;
aud[10536]=16'h3c3f;
aud[10537]=16'h3c46;
aud[10538]=16'h3c4d;
aud[10539]=16'h3c54;
aud[10540]=16'h3c5b;
aud[10541]=16'h3c63;
aud[10542]=16'h3c6a;
aud[10543]=16'h3c71;
aud[10544]=16'h3c78;
aud[10545]=16'h3c7f;
aud[10546]=16'h3c86;
aud[10547]=16'h3c8d;
aud[10548]=16'h3c94;
aud[10549]=16'h3c9b;
aud[10550]=16'h3ca1;
aud[10551]=16'h3ca8;
aud[10552]=16'h3caf;
aud[10553]=16'h3cb6;
aud[10554]=16'h3cbd;
aud[10555]=16'h3cc3;
aud[10556]=16'h3cca;
aud[10557]=16'h3cd1;
aud[10558]=16'h3cd7;
aud[10559]=16'h3cde;
aud[10560]=16'h3ce5;
aud[10561]=16'h3ceb;
aud[10562]=16'h3cf2;
aud[10563]=16'h3cf8;
aud[10564]=16'h3cff;
aud[10565]=16'h3d05;
aud[10566]=16'h3d0c;
aud[10567]=16'h3d12;
aud[10568]=16'h3d19;
aud[10569]=16'h3d1f;
aud[10570]=16'h3d25;
aud[10571]=16'h3d2c;
aud[10572]=16'h3d32;
aud[10573]=16'h3d38;
aud[10574]=16'h3d3f;
aud[10575]=16'h3d45;
aud[10576]=16'h3d4b;
aud[10577]=16'h3d51;
aud[10578]=16'h3d57;
aud[10579]=16'h3d5d;
aud[10580]=16'h3d63;
aud[10581]=16'h3d69;
aud[10582]=16'h3d6f;
aud[10583]=16'h3d75;
aud[10584]=16'h3d7b;
aud[10585]=16'h3d81;
aud[10586]=16'h3d87;
aud[10587]=16'h3d8d;
aud[10588]=16'h3d93;
aud[10589]=16'h3d99;
aud[10590]=16'h3d9f;
aud[10591]=16'h3da4;
aud[10592]=16'h3daa;
aud[10593]=16'h3db0;
aud[10594]=16'h3db6;
aud[10595]=16'h3dbb;
aud[10596]=16'h3dc1;
aud[10597]=16'h3dc7;
aud[10598]=16'h3dcc;
aud[10599]=16'h3dd2;
aud[10600]=16'h3dd7;
aud[10601]=16'h3ddd;
aud[10602]=16'h3de2;
aud[10603]=16'h3de8;
aud[10604]=16'h3ded;
aud[10605]=16'h3df3;
aud[10606]=16'h3df8;
aud[10607]=16'h3dfd;
aud[10608]=16'h3e03;
aud[10609]=16'h3e08;
aud[10610]=16'h3e0d;
aud[10611]=16'h3e12;
aud[10612]=16'h3e18;
aud[10613]=16'h3e1d;
aud[10614]=16'h3e22;
aud[10615]=16'h3e27;
aud[10616]=16'h3e2c;
aud[10617]=16'h3e31;
aud[10618]=16'h3e36;
aud[10619]=16'h3e3b;
aud[10620]=16'h3e40;
aud[10621]=16'h3e45;
aud[10622]=16'h3e4a;
aud[10623]=16'h3e4f;
aud[10624]=16'h3e54;
aud[10625]=16'h3e59;
aud[10626]=16'h3e5e;
aud[10627]=16'h3e62;
aud[10628]=16'h3e67;
aud[10629]=16'h3e6c;
aud[10630]=16'h3e71;
aud[10631]=16'h3e75;
aud[10632]=16'h3e7a;
aud[10633]=16'h3e7f;
aud[10634]=16'h3e83;
aud[10635]=16'h3e88;
aud[10636]=16'h3e8c;
aud[10637]=16'h3e91;
aud[10638]=16'h3e95;
aud[10639]=16'h3e9a;
aud[10640]=16'h3e9e;
aud[10641]=16'h3ea3;
aud[10642]=16'h3ea7;
aud[10643]=16'h3eac;
aud[10644]=16'h3eb0;
aud[10645]=16'h3eb4;
aud[10646]=16'h3eb9;
aud[10647]=16'h3ebd;
aud[10648]=16'h3ec1;
aud[10649]=16'h3ec5;
aud[10650]=16'h3ec9;
aud[10651]=16'h3ecd;
aud[10652]=16'h3ed2;
aud[10653]=16'h3ed6;
aud[10654]=16'h3eda;
aud[10655]=16'h3ede;
aud[10656]=16'h3ee2;
aud[10657]=16'h3ee6;
aud[10658]=16'h3eea;
aud[10659]=16'h3eee;
aud[10660]=16'h3ef2;
aud[10661]=16'h3ef5;
aud[10662]=16'h3ef9;
aud[10663]=16'h3efd;
aud[10664]=16'h3f01;
aud[10665]=16'h3f05;
aud[10666]=16'h3f08;
aud[10667]=16'h3f0c;
aud[10668]=16'h3f10;
aud[10669]=16'h3f13;
aud[10670]=16'h3f17;
aud[10671]=16'h3f1b;
aud[10672]=16'h3f1e;
aud[10673]=16'h3f22;
aud[10674]=16'h3f25;
aud[10675]=16'h3f29;
aud[10676]=16'h3f2c;
aud[10677]=16'h3f30;
aud[10678]=16'h3f33;
aud[10679]=16'h3f36;
aud[10680]=16'h3f3a;
aud[10681]=16'h3f3d;
aud[10682]=16'h3f40;
aud[10683]=16'h3f43;
aud[10684]=16'h3f47;
aud[10685]=16'h3f4a;
aud[10686]=16'h3f4d;
aud[10687]=16'h3f50;
aud[10688]=16'h3f53;
aud[10689]=16'h3f56;
aud[10690]=16'h3f5a;
aud[10691]=16'h3f5d;
aud[10692]=16'h3f60;
aud[10693]=16'h3f63;
aud[10694]=16'h3f65;
aud[10695]=16'h3f68;
aud[10696]=16'h3f6b;
aud[10697]=16'h3f6e;
aud[10698]=16'h3f71;
aud[10699]=16'h3f74;
aud[10700]=16'h3f77;
aud[10701]=16'h3f79;
aud[10702]=16'h3f7c;
aud[10703]=16'h3f7f;
aud[10704]=16'h3f81;
aud[10705]=16'h3f84;
aud[10706]=16'h3f87;
aud[10707]=16'h3f89;
aud[10708]=16'h3f8c;
aud[10709]=16'h3f8e;
aud[10710]=16'h3f91;
aud[10711]=16'h3f93;
aud[10712]=16'h3f96;
aud[10713]=16'h3f98;
aud[10714]=16'h3f9b;
aud[10715]=16'h3f9d;
aud[10716]=16'h3f9f;
aud[10717]=16'h3fa2;
aud[10718]=16'h3fa4;
aud[10719]=16'h3fa6;
aud[10720]=16'h3fa8;
aud[10721]=16'h3fab;
aud[10722]=16'h3fad;
aud[10723]=16'h3faf;
aud[10724]=16'h3fb1;
aud[10725]=16'h3fb3;
aud[10726]=16'h3fb5;
aud[10727]=16'h3fb7;
aud[10728]=16'h3fb9;
aud[10729]=16'h3fbb;
aud[10730]=16'h3fbd;
aud[10731]=16'h3fbf;
aud[10732]=16'h3fc1;
aud[10733]=16'h3fc3;
aud[10734]=16'h3fc5;
aud[10735]=16'h3fc7;
aud[10736]=16'h3fc8;
aud[10737]=16'h3fca;
aud[10738]=16'h3fcc;
aud[10739]=16'h3fcd;
aud[10740]=16'h3fcf;
aud[10741]=16'h3fd1;
aud[10742]=16'h3fd2;
aud[10743]=16'h3fd4;
aud[10744]=16'h3fd6;
aud[10745]=16'h3fd7;
aud[10746]=16'h3fd9;
aud[10747]=16'h3fda;
aud[10748]=16'h3fdc;
aud[10749]=16'h3fdd;
aud[10750]=16'h3fde;
aud[10751]=16'h3fe0;
aud[10752]=16'h3fe1;
aud[10753]=16'h3fe2;
aud[10754]=16'h3fe4;
aud[10755]=16'h3fe5;
aud[10756]=16'h3fe6;
aud[10757]=16'h3fe7;
aud[10758]=16'h3fe8;
aud[10759]=16'h3fea;
aud[10760]=16'h3feb;
aud[10761]=16'h3fec;
aud[10762]=16'h3fed;
aud[10763]=16'h3fee;
aud[10764]=16'h3fef;
aud[10765]=16'h3ff0;
aud[10766]=16'h3ff1;
aud[10767]=16'h3ff2;
aud[10768]=16'h3ff3;
aud[10769]=16'h3ff3;
aud[10770]=16'h3ff4;
aud[10771]=16'h3ff5;
aud[10772]=16'h3ff6;
aud[10773]=16'h3ff7;
aud[10774]=16'h3ff7;
aud[10775]=16'h3ff8;
aud[10776]=16'h3ff9;
aud[10777]=16'h3ff9;
aud[10778]=16'h3ffa;
aud[10779]=16'h3ffa;
aud[10780]=16'h3ffb;
aud[10781]=16'h3ffb;
aud[10782]=16'h3ffc;
aud[10783]=16'h3ffc;
aud[10784]=16'h3ffd;
aud[10785]=16'h3ffd;
aud[10786]=16'h3ffe;
aud[10787]=16'h3ffe;
aud[10788]=16'h3ffe;
aud[10789]=16'h3fff;
aud[10790]=16'h3fff;
aud[10791]=16'h3fff;
aud[10792]=16'h3fff;
aud[10793]=16'h3fff;
aud[10794]=16'h4000;
aud[10795]=16'h4000;
aud[10796]=16'h4000;
aud[10797]=16'h4000;
aud[10798]=16'h4000;
aud[10799]=16'h4000;
aud[10800]=16'h4000;
aud[10801]=16'h4000;
aud[10802]=16'h4000;
aud[10803]=16'h4000;
aud[10804]=16'h4000;
aud[10805]=16'h3fff;
aud[10806]=16'h3fff;
aud[10807]=16'h3fff;
aud[10808]=16'h3fff;
aud[10809]=16'h3fff;
aud[10810]=16'h3ffe;
aud[10811]=16'h3ffe;
aud[10812]=16'h3ffe;
aud[10813]=16'h3ffd;
aud[10814]=16'h3ffd;
aud[10815]=16'h3ffc;
aud[10816]=16'h3ffc;
aud[10817]=16'h3ffb;
aud[10818]=16'h3ffb;
aud[10819]=16'h3ffa;
aud[10820]=16'h3ffa;
aud[10821]=16'h3ff9;
aud[10822]=16'h3ff9;
aud[10823]=16'h3ff8;
aud[10824]=16'h3ff7;
aud[10825]=16'h3ff7;
aud[10826]=16'h3ff6;
aud[10827]=16'h3ff5;
aud[10828]=16'h3ff4;
aud[10829]=16'h3ff3;
aud[10830]=16'h3ff3;
aud[10831]=16'h3ff2;
aud[10832]=16'h3ff1;
aud[10833]=16'h3ff0;
aud[10834]=16'h3fef;
aud[10835]=16'h3fee;
aud[10836]=16'h3fed;
aud[10837]=16'h3fec;
aud[10838]=16'h3feb;
aud[10839]=16'h3fea;
aud[10840]=16'h3fe8;
aud[10841]=16'h3fe7;
aud[10842]=16'h3fe6;
aud[10843]=16'h3fe5;
aud[10844]=16'h3fe4;
aud[10845]=16'h3fe2;
aud[10846]=16'h3fe1;
aud[10847]=16'h3fe0;
aud[10848]=16'h3fde;
aud[10849]=16'h3fdd;
aud[10850]=16'h3fdc;
aud[10851]=16'h3fda;
aud[10852]=16'h3fd9;
aud[10853]=16'h3fd7;
aud[10854]=16'h3fd6;
aud[10855]=16'h3fd4;
aud[10856]=16'h3fd2;
aud[10857]=16'h3fd1;
aud[10858]=16'h3fcf;
aud[10859]=16'h3fcd;
aud[10860]=16'h3fcc;
aud[10861]=16'h3fca;
aud[10862]=16'h3fc8;
aud[10863]=16'h3fc7;
aud[10864]=16'h3fc5;
aud[10865]=16'h3fc3;
aud[10866]=16'h3fc1;
aud[10867]=16'h3fbf;
aud[10868]=16'h3fbd;
aud[10869]=16'h3fbb;
aud[10870]=16'h3fb9;
aud[10871]=16'h3fb7;
aud[10872]=16'h3fb5;
aud[10873]=16'h3fb3;
aud[10874]=16'h3fb1;
aud[10875]=16'h3faf;
aud[10876]=16'h3fad;
aud[10877]=16'h3fab;
aud[10878]=16'h3fa8;
aud[10879]=16'h3fa6;
aud[10880]=16'h3fa4;
aud[10881]=16'h3fa2;
aud[10882]=16'h3f9f;
aud[10883]=16'h3f9d;
aud[10884]=16'h3f9b;
aud[10885]=16'h3f98;
aud[10886]=16'h3f96;
aud[10887]=16'h3f93;
aud[10888]=16'h3f91;
aud[10889]=16'h3f8e;
aud[10890]=16'h3f8c;
aud[10891]=16'h3f89;
aud[10892]=16'h3f87;
aud[10893]=16'h3f84;
aud[10894]=16'h3f81;
aud[10895]=16'h3f7f;
aud[10896]=16'h3f7c;
aud[10897]=16'h3f79;
aud[10898]=16'h3f77;
aud[10899]=16'h3f74;
aud[10900]=16'h3f71;
aud[10901]=16'h3f6e;
aud[10902]=16'h3f6b;
aud[10903]=16'h3f68;
aud[10904]=16'h3f65;
aud[10905]=16'h3f63;
aud[10906]=16'h3f60;
aud[10907]=16'h3f5d;
aud[10908]=16'h3f5a;
aud[10909]=16'h3f56;
aud[10910]=16'h3f53;
aud[10911]=16'h3f50;
aud[10912]=16'h3f4d;
aud[10913]=16'h3f4a;
aud[10914]=16'h3f47;
aud[10915]=16'h3f43;
aud[10916]=16'h3f40;
aud[10917]=16'h3f3d;
aud[10918]=16'h3f3a;
aud[10919]=16'h3f36;
aud[10920]=16'h3f33;
aud[10921]=16'h3f30;
aud[10922]=16'h3f2c;
aud[10923]=16'h3f29;
aud[10924]=16'h3f25;
aud[10925]=16'h3f22;
aud[10926]=16'h3f1e;
aud[10927]=16'h3f1b;
aud[10928]=16'h3f17;
aud[10929]=16'h3f13;
aud[10930]=16'h3f10;
aud[10931]=16'h3f0c;
aud[10932]=16'h3f08;
aud[10933]=16'h3f05;
aud[10934]=16'h3f01;
aud[10935]=16'h3efd;
aud[10936]=16'h3ef9;
aud[10937]=16'h3ef5;
aud[10938]=16'h3ef2;
aud[10939]=16'h3eee;
aud[10940]=16'h3eea;
aud[10941]=16'h3ee6;
aud[10942]=16'h3ee2;
aud[10943]=16'h3ede;
aud[10944]=16'h3eda;
aud[10945]=16'h3ed6;
aud[10946]=16'h3ed2;
aud[10947]=16'h3ecd;
aud[10948]=16'h3ec9;
aud[10949]=16'h3ec5;
aud[10950]=16'h3ec1;
aud[10951]=16'h3ebd;
aud[10952]=16'h3eb9;
aud[10953]=16'h3eb4;
aud[10954]=16'h3eb0;
aud[10955]=16'h3eac;
aud[10956]=16'h3ea7;
aud[10957]=16'h3ea3;
aud[10958]=16'h3e9e;
aud[10959]=16'h3e9a;
aud[10960]=16'h3e95;
aud[10961]=16'h3e91;
aud[10962]=16'h3e8c;
aud[10963]=16'h3e88;
aud[10964]=16'h3e83;
aud[10965]=16'h3e7f;
aud[10966]=16'h3e7a;
aud[10967]=16'h3e75;
aud[10968]=16'h3e71;
aud[10969]=16'h3e6c;
aud[10970]=16'h3e67;
aud[10971]=16'h3e62;
aud[10972]=16'h3e5e;
aud[10973]=16'h3e59;
aud[10974]=16'h3e54;
aud[10975]=16'h3e4f;
aud[10976]=16'h3e4a;
aud[10977]=16'h3e45;
aud[10978]=16'h3e40;
aud[10979]=16'h3e3b;
aud[10980]=16'h3e36;
aud[10981]=16'h3e31;
aud[10982]=16'h3e2c;
aud[10983]=16'h3e27;
aud[10984]=16'h3e22;
aud[10985]=16'h3e1d;
aud[10986]=16'h3e18;
aud[10987]=16'h3e12;
aud[10988]=16'h3e0d;
aud[10989]=16'h3e08;
aud[10990]=16'h3e03;
aud[10991]=16'h3dfd;
aud[10992]=16'h3df8;
aud[10993]=16'h3df3;
aud[10994]=16'h3ded;
aud[10995]=16'h3de8;
aud[10996]=16'h3de2;
aud[10997]=16'h3ddd;
aud[10998]=16'h3dd7;
aud[10999]=16'h3dd2;
aud[11000]=16'h3dcc;
aud[11001]=16'h3dc7;
aud[11002]=16'h3dc1;
aud[11003]=16'h3dbb;
aud[11004]=16'h3db6;
aud[11005]=16'h3db0;
aud[11006]=16'h3daa;
aud[11007]=16'h3da4;
aud[11008]=16'h3d9f;
aud[11009]=16'h3d99;
aud[11010]=16'h3d93;
aud[11011]=16'h3d8d;
aud[11012]=16'h3d87;
aud[11013]=16'h3d81;
aud[11014]=16'h3d7b;
aud[11015]=16'h3d75;
aud[11016]=16'h3d6f;
aud[11017]=16'h3d69;
aud[11018]=16'h3d63;
aud[11019]=16'h3d5d;
aud[11020]=16'h3d57;
aud[11021]=16'h3d51;
aud[11022]=16'h3d4b;
aud[11023]=16'h3d45;
aud[11024]=16'h3d3f;
aud[11025]=16'h3d38;
aud[11026]=16'h3d32;
aud[11027]=16'h3d2c;
aud[11028]=16'h3d25;
aud[11029]=16'h3d1f;
aud[11030]=16'h3d19;
aud[11031]=16'h3d12;
aud[11032]=16'h3d0c;
aud[11033]=16'h3d05;
aud[11034]=16'h3cff;
aud[11035]=16'h3cf8;
aud[11036]=16'h3cf2;
aud[11037]=16'h3ceb;
aud[11038]=16'h3ce5;
aud[11039]=16'h3cde;
aud[11040]=16'h3cd7;
aud[11041]=16'h3cd1;
aud[11042]=16'h3cca;
aud[11043]=16'h3cc3;
aud[11044]=16'h3cbd;
aud[11045]=16'h3cb6;
aud[11046]=16'h3caf;
aud[11047]=16'h3ca8;
aud[11048]=16'h3ca1;
aud[11049]=16'h3c9b;
aud[11050]=16'h3c94;
aud[11051]=16'h3c8d;
aud[11052]=16'h3c86;
aud[11053]=16'h3c7f;
aud[11054]=16'h3c78;
aud[11055]=16'h3c71;
aud[11056]=16'h3c6a;
aud[11057]=16'h3c63;
aud[11058]=16'h3c5b;
aud[11059]=16'h3c54;
aud[11060]=16'h3c4d;
aud[11061]=16'h3c46;
aud[11062]=16'h3c3f;
aud[11063]=16'h3c37;
aud[11064]=16'h3c30;
aud[11065]=16'h3c29;
aud[11066]=16'h3c21;
aud[11067]=16'h3c1a;
aud[11068]=16'h3c13;
aud[11069]=16'h3c0b;
aud[11070]=16'h3c04;
aud[11071]=16'h3bfc;
aud[11072]=16'h3bf5;
aud[11073]=16'h3bed;
aud[11074]=16'h3be6;
aud[11075]=16'h3bde;
aud[11076]=16'h3bd7;
aud[11077]=16'h3bcf;
aud[11078]=16'h3bc7;
aud[11079]=16'h3bc0;
aud[11080]=16'h3bb8;
aud[11081]=16'h3bb0;
aud[11082]=16'h3ba9;
aud[11083]=16'h3ba1;
aud[11084]=16'h3b99;
aud[11085]=16'h3b91;
aud[11086]=16'h3b89;
aud[11087]=16'h3b81;
aud[11088]=16'h3b7a;
aud[11089]=16'h3b72;
aud[11090]=16'h3b6a;
aud[11091]=16'h3b62;
aud[11092]=16'h3b5a;
aud[11093]=16'h3b52;
aud[11094]=16'h3b4a;
aud[11095]=16'h3b41;
aud[11096]=16'h3b39;
aud[11097]=16'h3b31;
aud[11098]=16'h3b29;
aud[11099]=16'h3b21;
aud[11100]=16'h3b19;
aud[11101]=16'h3b10;
aud[11102]=16'h3b08;
aud[11103]=16'h3b00;
aud[11104]=16'h3af7;
aud[11105]=16'h3aef;
aud[11106]=16'h3ae7;
aud[11107]=16'h3ade;
aud[11108]=16'h3ad6;
aud[11109]=16'h3acd;
aud[11110]=16'h3ac5;
aud[11111]=16'h3abc;
aud[11112]=16'h3ab4;
aud[11113]=16'h3aab;
aud[11114]=16'h3aa3;
aud[11115]=16'h3a9a;
aud[11116]=16'h3a92;
aud[11117]=16'h3a89;
aud[11118]=16'h3a80;
aud[11119]=16'h3a78;
aud[11120]=16'h3a6f;
aud[11121]=16'h3a66;
aud[11122]=16'h3a5d;
aud[11123]=16'h3a54;
aud[11124]=16'h3a4c;
aud[11125]=16'h3a43;
aud[11126]=16'h3a3a;
aud[11127]=16'h3a31;
aud[11128]=16'h3a28;
aud[11129]=16'h3a1f;
aud[11130]=16'h3a16;
aud[11131]=16'h3a0d;
aud[11132]=16'h3a04;
aud[11133]=16'h39fb;
aud[11134]=16'h39f2;
aud[11135]=16'h39e9;
aud[11136]=16'h39e0;
aud[11137]=16'h39d6;
aud[11138]=16'h39cd;
aud[11139]=16'h39c4;
aud[11140]=16'h39bb;
aud[11141]=16'h39b1;
aud[11142]=16'h39a8;
aud[11143]=16'h399f;
aud[11144]=16'h3995;
aud[11145]=16'h398c;
aud[11146]=16'h3983;
aud[11147]=16'h3979;
aud[11148]=16'h3970;
aud[11149]=16'h3966;
aud[11150]=16'h395d;
aud[11151]=16'h3953;
aud[11152]=16'h394a;
aud[11153]=16'h3940;
aud[11154]=16'h3937;
aud[11155]=16'h392d;
aud[11156]=16'h3923;
aud[11157]=16'h391a;
aud[11158]=16'h3910;
aud[11159]=16'h3906;
aud[11160]=16'h38fd;
aud[11161]=16'h38f3;
aud[11162]=16'h38e9;
aud[11163]=16'h38df;
aud[11164]=16'h38d5;
aud[11165]=16'h38cb;
aud[11166]=16'h38c1;
aud[11167]=16'h38b8;
aud[11168]=16'h38ae;
aud[11169]=16'h38a4;
aud[11170]=16'h389a;
aud[11171]=16'h3890;
aud[11172]=16'h3886;
aud[11173]=16'h387b;
aud[11174]=16'h3871;
aud[11175]=16'h3867;
aud[11176]=16'h385d;
aud[11177]=16'h3853;
aud[11178]=16'h3849;
aud[11179]=16'h383f;
aud[11180]=16'h3834;
aud[11181]=16'h382a;
aud[11182]=16'h3820;
aud[11183]=16'h3815;
aud[11184]=16'h380b;
aud[11185]=16'h3801;
aud[11186]=16'h37f6;
aud[11187]=16'h37ec;
aud[11188]=16'h37e1;
aud[11189]=16'h37d7;
aud[11190]=16'h37cc;
aud[11191]=16'h37c2;
aud[11192]=16'h37b7;
aud[11193]=16'h37ad;
aud[11194]=16'h37a2;
aud[11195]=16'h3798;
aud[11196]=16'h378d;
aud[11197]=16'h3782;
aud[11198]=16'h3778;
aud[11199]=16'h376d;
aud[11200]=16'h3762;
aud[11201]=16'h3757;
aud[11202]=16'h374d;
aud[11203]=16'h3742;
aud[11204]=16'h3737;
aud[11205]=16'h372c;
aud[11206]=16'h3721;
aud[11207]=16'h3716;
aud[11208]=16'h370b;
aud[11209]=16'h3701;
aud[11210]=16'h36f6;
aud[11211]=16'h36eb;
aud[11212]=16'h36e0;
aud[11213]=16'h36d4;
aud[11214]=16'h36c9;
aud[11215]=16'h36be;
aud[11216]=16'h36b3;
aud[11217]=16'h36a8;
aud[11218]=16'h369d;
aud[11219]=16'h3692;
aud[11220]=16'h3686;
aud[11221]=16'h367b;
aud[11222]=16'h3670;
aud[11223]=16'h3665;
aud[11224]=16'h3659;
aud[11225]=16'h364e;
aud[11226]=16'h3643;
aud[11227]=16'h3637;
aud[11228]=16'h362c;
aud[11229]=16'h3620;
aud[11230]=16'h3615;
aud[11231]=16'h3609;
aud[11232]=16'h35fe;
aud[11233]=16'h35f2;
aud[11234]=16'h35e7;
aud[11235]=16'h35db;
aud[11236]=16'h35d0;
aud[11237]=16'h35c4;
aud[11238]=16'h35b8;
aud[11239]=16'h35ad;
aud[11240]=16'h35a1;
aud[11241]=16'h3595;
aud[11242]=16'h358a;
aud[11243]=16'h357e;
aud[11244]=16'h3572;
aud[11245]=16'h3566;
aud[11246]=16'h355a;
aud[11247]=16'h354f;
aud[11248]=16'h3543;
aud[11249]=16'h3537;
aud[11250]=16'h352b;
aud[11251]=16'h351f;
aud[11252]=16'h3513;
aud[11253]=16'h3507;
aud[11254]=16'h34fb;
aud[11255]=16'h34ef;
aud[11256]=16'h34e3;
aud[11257]=16'h34d7;
aud[11258]=16'h34cb;
aud[11259]=16'h34be;
aud[11260]=16'h34b2;
aud[11261]=16'h34a6;
aud[11262]=16'h349a;
aud[11263]=16'h348e;
aud[11264]=16'h3481;
aud[11265]=16'h3475;
aud[11266]=16'h3469;
aud[11267]=16'h345d;
aud[11268]=16'h3450;
aud[11269]=16'h3444;
aud[11270]=16'h3437;
aud[11271]=16'h342b;
aud[11272]=16'h341f;
aud[11273]=16'h3412;
aud[11274]=16'h3406;
aud[11275]=16'h33f9;
aud[11276]=16'h33ed;
aud[11277]=16'h33e0;
aud[11278]=16'h33d4;
aud[11279]=16'h33c7;
aud[11280]=16'h33ba;
aud[11281]=16'h33ae;
aud[11282]=16'h33a1;
aud[11283]=16'h3394;
aud[11284]=16'h3388;
aud[11285]=16'h337b;
aud[11286]=16'h336e;
aud[11287]=16'h3361;
aud[11288]=16'h3355;
aud[11289]=16'h3348;
aud[11290]=16'h333b;
aud[11291]=16'h332e;
aud[11292]=16'h3321;
aud[11293]=16'h3314;
aud[11294]=16'h3307;
aud[11295]=16'h32fa;
aud[11296]=16'h32ed;
aud[11297]=16'h32e0;
aud[11298]=16'h32d3;
aud[11299]=16'h32c6;
aud[11300]=16'h32b9;
aud[11301]=16'h32ac;
aud[11302]=16'h329f;
aud[11303]=16'h3292;
aud[11304]=16'h3285;
aud[11305]=16'h3278;
aud[11306]=16'h326a;
aud[11307]=16'h325d;
aud[11308]=16'h3250;
aud[11309]=16'h3243;
aud[11310]=16'h3235;
aud[11311]=16'h3228;
aud[11312]=16'h321b;
aud[11313]=16'h320d;
aud[11314]=16'h3200;
aud[11315]=16'h31f3;
aud[11316]=16'h31e5;
aud[11317]=16'h31d8;
aud[11318]=16'h31ca;
aud[11319]=16'h31bd;
aud[11320]=16'h31af;
aud[11321]=16'h31a2;
aud[11322]=16'h3194;
aud[11323]=16'h3187;
aud[11324]=16'h3179;
aud[11325]=16'h316b;
aud[11326]=16'h315e;
aud[11327]=16'h3150;
aud[11328]=16'h3142;
aud[11329]=16'h3135;
aud[11330]=16'h3127;
aud[11331]=16'h3119;
aud[11332]=16'h310b;
aud[11333]=16'h30fe;
aud[11334]=16'h30f0;
aud[11335]=16'h30e2;
aud[11336]=16'h30d4;
aud[11337]=16'h30c6;
aud[11338]=16'h30b8;
aud[11339]=16'h30aa;
aud[11340]=16'h309d;
aud[11341]=16'h308f;
aud[11342]=16'h3081;
aud[11343]=16'h3073;
aud[11344]=16'h3065;
aud[11345]=16'h3057;
aud[11346]=16'h3048;
aud[11347]=16'h303a;
aud[11348]=16'h302c;
aud[11349]=16'h301e;
aud[11350]=16'h3010;
aud[11351]=16'h3002;
aud[11352]=16'h2ff4;
aud[11353]=16'h2fe5;
aud[11354]=16'h2fd7;
aud[11355]=16'h2fc9;
aud[11356]=16'h2fbb;
aud[11357]=16'h2fac;
aud[11358]=16'h2f9e;
aud[11359]=16'h2f90;
aud[11360]=16'h2f81;
aud[11361]=16'h2f73;
aud[11362]=16'h2f65;
aud[11363]=16'h2f56;
aud[11364]=16'h2f48;
aud[11365]=16'h2f39;
aud[11366]=16'h2f2b;
aud[11367]=16'h2f1c;
aud[11368]=16'h2f0e;
aud[11369]=16'h2eff;
aud[11370]=16'h2ef1;
aud[11371]=16'h2ee2;
aud[11372]=16'h2ed3;
aud[11373]=16'h2ec5;
aud[11374]=16'h2eb6;
aud[11375]=16'h2ea7;
aud[11376]=16'h2e99;
aud[11377]=16'h2e8a;
aud[11378]=16'h2e7b;
aud[11379]=16'h2e6d;
aud[11380]=16'h2e5e;
aud[11381]=16'h2e4f;
aud[11382]=16'h2e40;
aud[11383]=16'h2e31;
aud[11384]=16'h2e22;
aud[11385]=16'h2e14;
aud[11386]=16'h2e05;
aud[11387]=16'h2df6;
aud[11388]=16'h2de7;
aud[11389]=16'h2dd8;
aud[11390]=16'h2dc9;
aud[11391]=16'h2dba;
aud[11392]=16'h2dab;
aud[11393]=16'h2d9c;
aud[11394]=16'h2d8d;
aud[11395]=16'h2d7e;
aud[11396]=16'h2d6f;
aud[11397]=16'h2d60;
aud[11398]=16'h2d50;
aud[11399]=16'h2d41;
aud[11400]=16'h2d32;
aud[11401]=16'h2d23;
aud[11402]=16'h2d14;
aud[11403]=16'h2d04;
aud[11404]=16'h2cf5;
aud[11405]=16'h2ce6;
aud[11406]=16'h2cd7;
aud[11407]=16'h2cc7;
aud[11408]=16'h2cb8;
aud[11409]=16'h2ca9;
aud[11410]=16'h2c99;
aud[11411]=16'h2c8a;
aud[11412]=16'h2c7a;
aud[11413]=16'h2c6b;
aud[11414]=16'h2c5c;
aud[11415]=16'h2c4c;
aud[11416]=16'h2c3d;
aud[11417]=16'h2c2d;
aud[11418]=16'h2c1e;
aud[11419]=16'h2c0e;
aud[11420]=16'h2bfe;
aud[11421]=16'h2bef;
aud[11422]=16'h2bdf;
aud[11423]=16'h2bd0;
aud[11424]=16'h2bc0;
aud[11425]=16'h2bb0;
aud[11426]=16'h2ba1;
aud[11427]=16'h2b91;
aud[11428]=16'h2b81;
aud[11429]=16'h2b71;
aud[11430]=16'h2b62;
aud[11431]=16'h2b52;
aud[11432]=16'h2b42;
aud[11433]=16'h2b32;
aud[11434]=16'h2b22;
aud[11435]=16'h2b13;
aud[11436]=16'h2b03;
aud[11437]=16'h2af3;
aud[11438]=16'h2ae3;
aud[11439]=16'h2ad3;
aud[11440]=16'h2ac3;
aud[11441]=16'h2ab3;
aud[11442]=16'h2aa3;
aud[11443]=16'h2a93;
aud[11444]=16'h2a83;
aud[11445]=16'h2a73;
aud[11446]=16'h2a63;
aud[11447]=16'h2a53;
aud[11448]=16'h2a43;
aud[11449]=16'h2a33;
aud[11450]=16'h2a23;
aud[11451]=16'h2a12;
aud[11452]=16'h2a02;
aud[11453]=16'h29f2;
aud[11454]=16'h29e2;
aud[11455]=16'h29d2;
aud[11456]=16'h29c1;
aud[11457]=16'h29b1;
aud[11458]=16'h29a1;
aud[11459]=16'h2991;
aud[11460]=16'h2980;
aud[11461]=16'h2970;
aud[11462]=16'h2960;
aud[11463]=16'h294f;
aud[11464]=16'h293f;
aud[11465]=16'h292e;
aud[11466]=16'h291e;
aud[11467]=16'h290e;
aud[11468]=16'h28fd;
aud[11469]=16'h28ed;
aud[11470]=16'h28dc;
aud[11471]=16'h28cc;
aud[11472]=16'h28bb;
aud[11473]=16'h28aa;
aud[11474]=16'h289a;
aud[11475]=16'h2889;
aud[11476]=16'h2879;
aud[11477]=16'h2868;
aud[11478]=16'h2857;
aud[11479]=16'h2847;
aud[11480]=16'h2836;
aud[11481]=16'h2825;
aud[11482]=16'h2815;
aud[11483]=16'h2804;
aud[11484]=16'h27f3;
aud[11485]=16'h27e2;
aud[11486]=16'h27d2;
aud[11487]=16'h27c1;
aud[11488]=16'h27b0;
aud[11489]=16'h279f;
aud[11490]=16'h278e;
aud[11491]=16'h277e;
aud[11492]=16'h276d;
aud[11493]=16'h275c;
aud[11494]=16'h274b;
aud[11495]=16'h273a;
aud[11496]=16'h2729;
aud[11497]=16'h2718;
aud[11498]=16'h2707;
aud[11499]=16'h26f6;
aud[11500]=16'h26e5;
aud[11501]=16'h26d4;
aud[11502]=16'h26c3;
aud[11503]=16'h26b2;
aud[11504]=16'h26a1;
aud[11505]=16'h2690;
aud[11506]=16'h267e;
aud[11507]=16'h266d;
aud[11508]=16'h265c;
aud[11509]=16'h264b;
aud[11510]=16'h263a;
aud[11511]=16'h2629;
aud[11512]=16'h2617;
aud[11513]=16'h2606;
aud[11514]=16'h25f5;
aud[11515]=16'h25e4;
aud[11516]=16'h25d2;
aud[11517]=16'h25c1;
aud[11518]=16'h25b0;
aud[11519]=16'h259e;
aud[11520]=16'h258d;
aud[11521]=16'h257c;
aud[11522]=16'h256a;
aud[11523]=16'h2559;
aud[11524]=16'h2547;
aud[11525]=16'h2536;
aud[11526]=16'h2524;
aud[11527]=16'h2513;
aud[11528]=16'h2501;
aud[11529]=16'h24f0;
aud[11530]=16'h24de;
aud[11531]=16'h24cd;
aud[11532]=16'h24bb;
aud[11533]=16'h24aa;
aud[11534]=16'h2498;
aud[11535]=16'h2487;
aud[11536]=16'h2475;
aud[11537]=16'h2463;
aud[11538]=16'h2452;
aud[11539]=16'h2440;
aud[11540]=16'h242e;
aud[11541]=16'h241d;
aud[11542]=16'h240b;
aud[11543]=16'h23f9;
aud[11544]=16'h23e7;
aud[11545]=16'h23d6;
aud[11546]=16'h23c4;
aud[11547]=16'h23b2;
aud[11548]=16'h23a0;
aud[11549]=16'h238e;
aud[11550]=16'h237d;
aud[11551]=16'h236b;
aud[11552]=16'h2359;
aud[11553]=16'h2347;
aud[11554]=16'h2335;
aud[11555]=16'h2323;
aud[11556]=16'h2311;
aud[11557]=16'h22ff;
aud[11558]=16'h22ed;
aud[11559]=16'h22db;
aud[11560]=16'h22c9;
aud[11561]=16'h22b7;
aud[11562]=16'h22a5;
aud[11563]=16'h2293;
aud[11564]=16'h2281;
aud[11565]=16'h226f;
aud[11566]=16'h225d;
aud[11567]=16'h224b;
aud[11568]=16'h2239;
aud[11569]=16'h2227;
aud[11570]=16'h2215;
aud[11571]=16'h2202;
aud[11572]=16'h21f0;
aud[11573]=16'h21de;
aud[11574]=16'h21cc;
aud[11575]=16'h21ba;
aud[11576]=16'h21a7;
aud[11577]=16'h2195;
aud[11578]=16'h2183;
aud[11579]=16'h2171;
aud[11580]=16'h215e;
aud[11581]=16'h214c;
aud[11582]=16'h213a;
aud[11583]=16'h2127;
aud[11584]=16'h2115;
aud[11585]=16'h2103;
aud[11586]=16'h20f0;
aud[11587]=16'h20de;
aud[11588]=16'h20cb;
aud[11589]=16'h20b9;
aud[11590]=16'h20a7;
aud[11591]=16'h2094;
aud[11592]=16'h2082;
aud[11593]=16'h206f;
aud[11594]=16'h205d;
aud[11595]=16'h204a;
aud[11596]=16'h2038;
aud[11597]=16'h2025;
aud[11598]=16'h2013;
aud[11599]=16'h2000;
aud[11600]=16'h1fed;
aud[11601]=16'h1fdb;
aud[11602]=16'h1fc8;
aud[11603]=16'h1fb6;
aud[11604]=16'h1fa3;
aud[11605]=16'h1f90;
aud[11606]=16'h1f7e;
aud[11607]=16'h1f6b;
aud[11608]=16'h1f58;
aud[11609]=16'h1f46;
aud[11610]=16'h1f33;
aud[11611]=16'h1f20;
aud[11612]=16'h1f0d;
aud[11613]=16'h1efb;
aud[11614]=16'h1ee8;
aud[11615]=16'h1ed5;
aud[11616]=16'h1ec2;
aud[11617]=16'h1eaf;
aud[11618]=16'h1e9d;
aud[11619]=16'h1e8a;
aud[11620]=16'h1e77;
aud[11621]=16'h1e64;
aud[11622]=16'h1e51;
aud[11623]=16'h1e3e;
aud[11624]=16'h1e2b;
aud[11625]=16'h1e18;
aud[11626]=16'h1e06;
aud[11627]=16'h1df3;
aud[11628]=16'h1de0;
aud[11629]=16'h1dcd;
aud[11630]=16'h1dba;
aud[11631]=16'h1da7;
aud[11632]=16'h1d94;
aud[11633]=16'h1d81;
aud[11634]=16'h1d6e;
aud[11635]=16'h1d5b;
aud[11636]=16'h1d47;
aud[11637]=16'h1d34;
aud[11638]=16'h1d21;
aud[11639]=16'h1d0e;
aud[11640]=16'h1cfb;
aud[11641]=16'h1ce8;
aud[11642]=16'h1cd5;
aud[11643]=16'h1cc2;
aud[11644]=16'h1cae;
aud[11645]=16'h1c9b;
aud[11646]=16'h1c88;
aud[11647]=16'h1c75;
aud[11648]=16'h1c62;
aud[11649]=16'h1c4e;
aud[11650]=16'h1c3b;
aud[11651]=16'h1c28;
aud[11652]=16'h1c15;
aud[11653]=16'h1c01;
aud[11654]=16'h1bee;
aud[11655]=16'h1bdb;
aud[11656]=16'h1bc8;
aud[11657]=16'h1bb4;
aud[11658]=16'h1ba1;
aud[11659]=16'h1b8d;
aud[11660]=16'h1b7a;
aud[11661]=16'h1b67;
aud[11662]=16'h1b53;
aud[11663]=16'h1b40;
aud[11664]=16'h1b2d;
aud[11665]=16'h1b19;
aud[11666]=16'h1b06;
aud[11667]=16'h1af2;
aud[11668]=16'h1adf;
aud[11669]=16'h1acb;
aud[11670]=16'h1ab8;
aud[11671]=16'h1aa4;
aud[11672]=16'h1a91;
aud[11673]=16'h1a7d;
aud[11674]=16'h1a6a;
aud[11675]=16'h1a56;
aud[11676]=16'h1a43;
aud[11677]=16'h1a2f;
aud[11678]=16'h1a1c;
aud[11679]=16'h1a08;
aud[11680]=16'h19f4;
aud[11681]=16'h19e1;
aud[11682]=16'h19cd;
aud[11683]=16'h19ba;
aud[11684]=16'h19a6;
aud[11685]=16'h1992;
aud[11686]=16'h197f;
aud[11687]=16'h196b;
aud[11688]=16'h1957;
aud[11689]=16'h1943;
aud[11690]=16'h1930;
aud[11691]=16'h191c;
aud[11692]=16'h1908;
aud[11693]=16'h18f5;
aud[11694]=16'h18e1;
aud[11695]=16'h18cd;
aud[11696]=16'h18b9;
aud[11697]=16'h18a5;
aud[11698]=16'h1892;
aud[11699]=16'h187e;
aud[11700]=16'h186a;
aud[11701]=16'h1856;
aud[11702]=16'h1842;
aud[11703]=16'h182f;
aud[11704]=16'h181b;
aud[11705]=16'h1807;
aud[11706]=16'h17f3;
aud[11707]=16'h17df;
aud[11708]=16'h17cb;
aud[11709]=16'h17b7;
aud[11710]=16'h17a3;
aud[11711]=16'h178f;
aud[11712]=16'h177b;
aud[11713]=16'h1767;
aud[11714]=16'h1753;
aud[11715]=16'h1740;
aud[11716]=16'h172c;
aud[11717]=16'h1718;
aud[11718]=16'h1704;
aud[11719]=16'h16f0;
aud[11720]=16'h16db;
aud[11721]=16'h16c7;
aud[11722]=16'h16b3;
aud[11723]=16'h169f;
aud[11724]=16'h168b;
aud[11725]=16'h1677;
aud[11726]=16'h1663;
aud[11727]=16'h164f;
aud[11728]=16'h163b;
aud[11729]=16'h1627;
aud[11730]=16'h1613;
aud[11731]=16'h15ff;
aud[11732]=16'h15ea;
aud[11733]=16'h15d6;
aud[11734]=16'h15c2;
aud[11735]=16'h15ae;
aud[11736]=16'h159a;
aud[11737]=16'h1586;
aud[11738]=16'h1571;
aud[11739]=16'h155d;
aud[11740]=16'h1549;
aud[11741]=16'h1535;
aud[11742]=16'h1520;
aud[11743]=16'h150c;
aud[11744]=16'h14f8;
aud[11745]=16'h14e4;
aud[11746]=16'h14cf;
aud[11747]=16'h14bb;
aud[11748]=16'h14a7;
aud[11749]=16'h1492;
aud[11750]=16'h147e;
aud[11751]=16'h146a;
aud[11752]=16'h1455;
aud[11753]=16'h1441;
aud[11754]=16'h142d;
aud[11755]=16'h1418;
aud[11756]=16'h1404;
aud[11757]=16'h13f0;
aud[11758]=16'h13db;
aud[11759]=16'h13c7;
aud[11760]=16'h13b3;
aud[11761]=16'h139e;
aud[11762]=16'h138a;
aud[11763]=16'h1375;
aud[11764]=16'h1361;
aud[11765]=16'h134c;
aud[11766]=16'h1338;
aud[11767]=16'h1323;
aud[11768]=16'h130f;
aud[11769]=16'h12fb;
aud[11770]=16'h12e6;
aud[11771]=16'h12d2;
aud[11772]=16'h12bd;
aud[11773]=16'h12a9;
aud[11774]=16'h1294;
aud[11775]=16'h127f;
aud[11776]=16'h126b;
aud[11777]=16'h1256;
aud[11778]=16'h1242;
aud[11779]=16'h122d;
aud[11780]=16'h1219;
aud[11781]=16'h1204;
aud[11782]=16'h11f0;
aud[11783]=16'h11db;
aud[11784]=16'h11c6;
aud[11785]=16'h11b2;
aud[11786]=16'h119d;
aud[11787]=16'h1189;
aud[11788]=16'h1174;
aud[11789]=16'h115f;
aud[11790]=16'h114b;
aud[11791]=16'h1136;
aud[11792]=16'h1121;
aud[11793]=16'h110d;
aud[11794]=16'h10f8;
aud[11795]=16'h10e3;
aud[11796]=16'h10cf;
aud[11797]=16'h10ba;
aud[11798]=16'h10a5;
aud[11799]=16'h1090;
aud[11800]=16'h107c;
aud[11801]=16'h1067;
aud[11802]=16'h1052;
aud[11803]=16'h103e;
aud[11804]=16'h1029;
aud[11805]=16'h1014;
aud[11806]=16'hfff;
aud[11807]=16'hfeb;
aud[11808]=16'hfd6;
aud[11809]=16'hfc1;
aud[11810]=16'hfac;
aud[11811]=16'hf97;
aud[11812]=16'hf83;
aud[11813]=16'hf6e;
aud[11814]=16'hf59;
aud[11815]=16'hf44;
aud[11816]=16'hf2f;
aud[11817]=16'hf1a;
aud[11818]=16'hf06;
aud[11819]=16'hef1;
aud[11820]=16'hedc;
aud[11821]=16'hec7;
aud[11822]=16'heb2;
aud[11823]=16'he9d;
aud[11824]=16'he88;
aud[11825]=16'he74;
aud[11826]=16'he5f;
aud[11827]=16'he4a;
aud[11828]=16'he35;
aud[11829]=16'he20;
aud[11830]=16'he0b;
aud[11831]=16'hdf6;
aud[11832]=16'hde1;
aud[11833]=16'hdcc;
aud[11834]=16'hdb7;
aud[11835]=16'hda2;
aud[11836]=16'hd8d;
aud[11837]=16'hd78;
aud[11838]=16'hd63;
aud[11839]=16'hd4e;
aud[11840]=16'hd39;
aud[11841]=16'hd24;
aud[11842]=16'hd0f;
aud[11843]=16'hcfa;
aud[11844]=16'hce5;
aud[11845]=16'hcd0;
aud[11846]=16'hcbb;
aud[11847]=16'hca6;
aud[11848]=16'hc91;
aud[11849]=16'hc7c;
aud[11850]=16'hc67;
aud[11851]=16'hc52;
aud[11852]=16'hc3d;
aud[11853]=16'hc28;
aud[11854]=16'hc13;
aud[11855]=16'hbfe;
aud[11856]=16'hbe9;
aud[11857]=16'hbd4;
aud[11858]=16'hbbf;
aud[11859]=16'hbaa;
aud[11860]=16'hb95;
aud[11861]=16'hb80;
aud[11862]=16'hb6a;
aud[11863]=16'hb55;
aud[11864]=16'hb40;
aud[11865]=16'hb2b;
aud[11866]=16'hb16;
aud[11867]=16'hb01;
aud[11868]=16'haec;
aud[11869]=16'had7;
aud[11870]=16'hac1;
aud[11871]=16'haac;
aud[11872]=16'ha97;
aud[11873]=16'ha82;
aud[11874]=16'ha6d;
aud[11875]=16'ha58;
aud[11876]=16'ha43;
aud[11877]=16'ha2d;
aud[11878]=16'ha18;
aud[11879]=16'ha03;
aud[11880]=16'h9ee;
aud[11881]=16'h9d9;
aud[11882]=16'h9c3;
aud[11883]=16'h9ae;
aud[11884]=16'h999;
aud[11885]=16'h984;
aud[11886]=16'h96f;
aud[11887]=16'h959;
aud[11888]=16'h944;
aud[11889]=16'h92f;
aud[11890]=16'h91a;
aud[11891]=16'h905;
aud[11892]=16'h8ef;
aud[11893]=16'h8da;
aud[11894]=16'h8c5;
aud[11895]=16'h8b0;
aud[11896]=16'h89a;
aud[11897]=16'h885;
aud[11898]=16'h870;
aud[11899]=16'h85b;
aud[11900]=16'h845;
aud[11901]=16'h830;
aud[11902]=16'h81b;
aud[11903]=16'h805;
aud[11904]=16'h7f0;
aud[11905]=16'h7db;
aud[11906]=16'h7c6;
aud[11907]=16'h7b0;
aud[11908]=16'h79b;
aud[11909]=16'h786;
aud[11910]=16'h770;
aud[11911]=16'h75b;
aud[11912]=16'h746;
aud[11913]=16'h731;
aud[11914]=16'h71b;
aud[11915]=16'h706;
aud[11916]=16'h6f1;
aud[11917]=16'h6db;
aud[11918]=16'h6c6;
aud[11919]=16'h6b1;
aud[11920]=16'h69b;
aud[11921]=16'h686;
aud[11922]=16'h671;
aud[11923]=16'h65b;
aud[11924]=16'h646;
aud[11925]=16'h631;
aud[11926]=16'h61b;
aud[11927]=16'h606;
aud[11928]=16'h5f1;
aud[11929]=16'h5db;
aud[11930]=16'h5c6;
aud[11931]=16'h5b0;
aud[11932]=16'h59b;
aud[11933]=16'h586;
aud[11934]=16'h570;
aud[11935]=16'h55b;
aud[11936]=16'h546;
aud[11937]=16'h530;
aud[11938]=16'h51b;
aud[11939]=16'h505;
aud[11940]=16'h4f0;
aud[11941]=16'h4db;
aud[11942]=16'h4c5;
aud[11943]=16'h4b0;
aud[11944]=16'h49b;
aud[11945]=16'h485;
aud[11946]=16'h470;
aud[11947]=16'h45a;
aud[11948]=16'h445;
aud[11949]=16'h430;
aud[11950]=16'h41a;
aud[11951]=16'h405;
aud[11952]=16'h3ef;
aud[11953]=16'h3da;
aud[11954]=16'h3c5;
aud[11955]=16'h3af;
aud[11956]=16'h39a;
aud[11957]=16'h384;
aud[11958]=16'h36f;
aud[11959]=16'h359;
aud[11960]=16'h344;
aud[11961]=16'h32f;
aud[11962]=16'h319;
aud[11963]=16'h304;
aud[11964]=16'h2ee;
aud[11965]=16'h2d9;
aud[11966]=16'h2c4;
aud[11967]=16'h2ae;
aud[11968]=16'h299;
aud[11969]=16'h283;
aud[11970]=16'h26e;
aud[11971]=16'h258;
aud[11972]=16'h243;
aud[11973]=16'h22e;
aud[11974]=16'h218;
aud[11975]=16'h203;
aud[11976]=16'h1ed;
aud[11977]=16'h1d8;
aud[11978]=16'h1c2;
aud[11979]=16'h1ad;
aud[11980]=16'h197;
aud[11981]=16'h182;
aud[11982]=16'h16d;
aud[11983]=16'h157;
aud[11984]=16'h142;
aud[11985]=16'h12c;
aud[11986]=16'h117;
aud[11987]=16'h101;
aud[11988]=16'hec;
aud[11989]=16'hd6;
aud[11990]=16'hc1;
aud[11991]=16'hac;
aud[11992]=16'h96;
aud[11993]=16'h81;
aud[11994]=16'h6b;
aud[11995]=16'h56;
aud[11996]=16'h40;
aud[11997]=16'h2b;
aud[11998]=16'h15;
aud[11999]=16'h0;
aud[12000]=16'hffeb;
aud[12001]=16'hffd5;
aud[12002]=16'hffc0;
aud[12003]=16'hffaa;
aud[12004]=16'hff95;
aud[12005]=16'hff7f;
aud[12006]=16'hff6a;
aud[12007]=16'hff54;
aud[12008]=16'hff3f;
aud[12009]=16'hff2a;
aud[12010]=16'hff14;
aud[12011]=16'hfeff;
aud[12012]=16'hfee9;
aud[12013]=16'hfed4;
aud[12014]=16'hfebe;
aud[12015]=16'hfea9;
aud[12016]=16'hfe93;
aud[12017]=16'hfe7e;
aud[12018]=16'hfe69;
aud[12019]=16'hfe53;
aud[12020]=16'hfe3e;
aud[12021]=16'hfe28;
aud[12022]=16'hfe13;
aud[12023]=16'hfdfd;
aud[12024]=16'hfde8;
aud[12025]=16'hfdd2;
aud[12026]=16'hfdbd;
aud[12027]=16'hfda8;
aud[12028]=16'hfd92;
aud[12029]=16'hfd7d;
aud[12030]=16'hfd67;
aud[12031]=16'hfd52;
aud[12032]=16'hfd3c;
aud[12033]=16'hfd27;
aud[12034]=16'hfd12;
aud[12035]=16'hfcfc;
aud[12036]=16'hfce7;
aud[12037]=16'hfcd1;
aud[12038]=16'hfcbc;
aud[12039]=16'hfca7;
aud[12040]=16'hfc91;
aud[12041]=16'hfc7c;
aud[12042]=16'hfc66;
aud[12043]=16'hfc51;
aud[12044]=16'hfc3b;
aud[12045]=16'hfc26;
aud[12046]=16'hfc11;
aud[12047]=16'hfbfb;
aud[12048]=16'hfbe6;
aud[12049]=16'hfbd0;
aud[12050]=16'hfbbb;
aud[12051]=16'hfba6;
aud[12052]=16'hfb90;
aud[12053]=16'hfb7b;
aud[12054]=16'hfb65;
aud[12055]=16'hfb50;
aud[12056]=16'hfb3b;
aud[12057]=16'hfb25;
aud[12058]=16'hfb10;
aud[12059]=16'hfafb;
aud[12060]=16'hfae5;
aud[12061]=16'hfad0;
aud[12062]=16'hfaba;
aud[12063]=16'hfaa5;
aud[12064]=16'hfa90;
aud[12065]=16'hfa7a;
aud[12066]=16'hfa65;
aud[12067]=16'hfa50;
aud[12068]=16'hfa3a;
aud[12069]=16'hfa25;
aud[12070]=16'hfa0f;
aud[12071]=16'hf9fa;
aud[12072]=16'hf9e5;
aud[12073]=16'hf9cf;
aud[12074]=16'hf9ba;
aud[12075]=16'hf9a5;
aud[12076]=16'hf98f;
aud[12077]=16'hf97a;
aud[12078]=16'hf965;
aud[12079]=16'hf94f;
aud[12080]=16'hf93a;
aud[12081]=16'hf925;
aud[12082]=16'hf90f;
aud[12083]=16'hf8fa;
aud[12084]=16'hf8e5;
aud[12085]=16'hf8cf;
aud[12086]=16'hf8ba;
aud[12087]=16'hf8a5;
aud[12088]=16'hf890;
aud[12089]=16'hf87a;
aud[12090]=16'hf865;
aud[12091]=16'hf850;
aud[12092]=16'hf83a;
aud[12093]=16'hf825;
aud[12094]=16'hf810;
aud[12095]=16'hf7fb;
aud[12096]=16'hf7e5;
aud[12097]=16'hf7d0;
aud[12098]=16'hf7bb;
aud[12099]=16'hf7a5;
aud[12100]=16'hf790;
aud[12101]=16'hf77b;
aud[12102]=16'hf766;
aud[12103]=16'hf750;
aud[12104]=16'hf73b;
aud[12105]=16'hf726;
aud[12106]=16'hf711;
aud[12107]=16'hf6fb;
aud[12108]=16'hf6e6;
aud[12109]=16'hf6d1;
aud[12110]=16'hf6bc;
aud[12111]=16'hf6a7;
aud[12112]=16'hf691;
aud[12113]=16'hf67c;
aud[12114]=16'hf667;
aud[12115]=16'hf652;
aud[12116]=16'hf63d;
aud[12117]=16'hf627;
aud[12118]=16'hf612;
aud[12119]=16'hf5fd;
aud[12120]=16'hf5e8;
aud[12121]=16'hf5d3;
aud[12122]=16'hf5bd;
aud[12123]=16'hf5a8;
aud[12124]=16'hf593;
aud[12125]=16'hf57e;
aud[12126]=16'hf569;
aud[12127]=16'hf554;
aud[12128]=16'hf53f;
aud[12129]=16'hf529;
aud[12130]=16'hf514;
aud[12131]=16'hf4ff;
aud[12132]=16'hf4ea;
aud[12133]=16'hf4d5;
aud[12134]=16'hf4c0;
aud[12135]=16'hf4ab;
aud[12136]=16'hf496;
aud[12137]=16'hf480;
aud[12138]=16'hf46b;
aud[12139]=16'hf456;
aud[12140]=16'hf441;
aud[12141]=16'hf42c;
aud[12142]=16'hf417;
aud[12143]=16'hf402;
aud[12144]=16'hf3ed;
aud[12145]=16'hf3d8;
aud[12146]=16'hf3c3;
aud[12147]=16'hf3ae;
aud[12148]=16'hf399;
aud[12149]=16'hf384;
aud[12150]=16'hf36f;
aud[12151]=16'hf35a;
aud[12152]=16'hf345;
aud[12153]=16'hf330;
aud[12154]=16'hf31b;
aud[12155]=16'hf306;
aud[12156]=16'hf2f1;
aud[12157]=16'hf2dc;
aud[12158]=16'hf2c7;
aud[12159]=16'hf2b2;
aud[12160]=16'hf29d;
aud[12161]=16'hf288;
aud[12162]=16'hf273;
aud[12163]=16'hf25e;
aud[12164]=16'hf249;
aud[12165]=16'hf234;
aud[12166]=16'hf21f;
aud[12167]=16'hf20a;
aud[12168]=16'hf1f5;
aud[12169]=16'hf1e0;
aud[12170]=16'hf1cb;
aud[12171]=16'hf1b6;
aud[12172]=16'hf1a1;
aud[12173]=16'hf18c;
aud[12174]=16'hf178;
aud[12175]=16'hf163;
aud[12176]=16'hf14e;
aud[12177]=16'hf139;
aud[12178]=16'hf124;
aud[12179]=16'hf10f;
aud[12180]=16'hf0fa;
aud[12181]=16'hf0e6;
aud[12182]=16'hf0d1;
aud[12183]=16'hf0bc;
aud[12184]=16'hf0a7;
aud[12185]=16'hf092;
aud[12186]=16'hf07d;
aud[12187]=16'hf069;
aud[12188]=16'hf054;
aud[12189]=16'hf03f;
aud[12190]=16'hf02a;
aud[12191]=16'hf015;
aud[12192]=16'hf001;
aud[12193]=16'hefec;
aud[12194]=16'hefd7;
aud[12195]=16'hefc2;
aud[12196]=16'hefae;
aud[12197]=16'hef99;
aud[12198]=16'hef84;
aud[12199]=16'hef70;
aud[12200]=16'hef5b;
aud[12201]=16'hef46;
aud[12202]=16'hef31;
aud[12203]=16'hef1d;
aud[12204]=16'hef08;
aud[12205]=16'heef3;
aud[12206]=16'heedf;
aud[12207]=16'heeca;
aud[12208]=16'heeb5;
aud[12209]=16'heea1;
aud[12210]=16'hee8c;
aud[12211]=16'hee77;
aud[12212]=16'hee63;
aud[12213]=16'hee4e;
aud[12214]=16'hee3a;
aud[12215]=16'hee25;
aud[12216]=16'hee10;
aud[12217]=16'hedfc;
aud[12218]=16'hede7;
aud[12219]=16'hedd3;
aud[12220]=16'hedbe;
aud[12221]=16'hedaa;
aud[12222]=16'hed95;
aud[12223]=16'hed81;
aud[12224]=16'hed6c;
aud[12225]=16'hed57;
aud[12226]=16'hed43;
aud[12227]=16'hed2e;
aud[12228]=16'hed1a;
aud[12229]=16'hed05;
aud[12230]=16'hecf1;
aud[12231]=16'hecdd;
aud[12232]=16'hecc8;
aud[12233]=16'hecb4;
aud[12234]=16'hec9f;
aud[12235]=16'hec8b;
aud[12236]=16'hec76;
aud[12237]=16'hec62;
aud[12238]=16'hec4d;
aud[12239]=16'hec39;
aud[12240]=16'hec25;
aud[12241]=16'hec10;
aud[12242]=16'hebfc;
aud[12243]=16'hebe8;
aud[12244]=16'hebd3;
aud[12245]=16'hebbf;
aud[12246]=16'hebab;
aud[12247]=16'heb96;
aud[12248]=16'heb82;
aud[12249]=16'heb6e;
aud[12250]=16'heb59;
aud[12251]=16'heb45;
aud[12252]=16'heb31;
aud[12253]=16'heb1c;
aud[12254]=16'heb08;
aud[12255]=16'heaf4;
aud[12256]=16'heae0;
aud[12257]=16'heacb;
aud[12258]=16'heab7;
aud[12259]=16'heaa3;
aud[12260]=16'hea8f;
aud[12261]=16'hea7a;
aud[12262]=16'hea66;
aud[12263]=16'hea52;
aud[12264]=16'hea3e;
aud[12265]=16'hea2a;
aud[12266]=16'hea16;
aud[12267]=16'hea01;
aud[12268]=16'he9ed;
aud[12269]=16'he9d9;
aud[12270]=16'he9c5;
aud[12271]=16'he9b1;
aud[12272]=16'he99d;
aud[12273]=16'he989;
aud[12274]=16'he975;
aud[12275]=16'he961;
aud[12276]=16'he94d;
aud[12277]=16'he939;
aud[12278]=16'he925;
aud[12279]=16'he910;
aud[12280]=16'he8fc;
aud[12281]=16'he8e8;
aud[12282]=16'he8d4;
aud[12283]=16'he8c0;
aud[12284]=16'he8ad;
aud[12285]=16'he899;
aud[12286]=16'he885;
aud[12287]=16'he871;
aud[12288]=16'he85d;
aud[12289]=16'he849;
aud[12290]=16'he835;
aud[12291]=16'he821;
aud[12292]=16'he80d;
aud[12293]=16'he7f9;
aud[12294]=16'he7e5;
aud[12295]=16'he7d1;
aud[12296]=16'he7be;
aud[12297]=16'he7aa;
aud[12298]=16'he796;
aud[12299]=16'he782;
aud[12300]=16'he76e;
aud[12301]=16'he75b;
aud[12302]=16'he747;
aud[12303]=16'he733;
aud[12304]=16'he71f;
aud[12305]=16'he70b;
aud[12306]=16'he6f8;
aud[12307]=16'he6e4;
aud[12308]=16'he6d0;
aud[12309]=16'he6bd;
aud[12310]=16'he6a9;
aud[12311]=16'he695;
aud[12312]=16'he681;
aud[12313]=16'he66e;
aud[12314]=16'he65a;
aud[12315]=16'he646;
aud[12316]=16'he633;
aud[12317]=16'he61f;
aud[12318]=16'he60c;
aud[12319]=16'he5f8;
aud[12320]=16'he5e4;
aud[12321]=16'he5d1;
aud[12322]=16'he5bd;
aud[12323]=16'he5aa;
aud[12324]=16'he596;
aud[12325]=16'he583;
aud[12326]=16'he56f;
aud[12327]=16'he55c;
aud[12328]=16'he548;
aud[12329]=16'he535;
aud[12330]=16'he521;
aud[12331]=16'he50e;
aud[12332]=16'he4fa;
aud[12333]=16'he4e7;
aud[12334]=16'he4d3;
aud[12335]=16'he4c0;
aud[12336]=16'he4ad;
aud[12337]=16'he499;
aud[12338]=16'he486;
aud[12339]=16'he473;
aud[12340]=16'he45f;
aud[12341]=16'he44c;
aud[12342]=16'he438;
aud[12343]=16'he425;
aud[12344]=16'he412;
aud[12345]=16'he3ff;
aud[12346]=16'he3eb;
aud[12347]=16'he3d8;
aud[12348]=16'he3c5;
aud[12349]=16'he3b2;
aud[12350]=16'he39e;
aud[12351]=16'he38b;
aud[12352]=16'he378;
aud[12353]=16'he365;
aud[12354]=16'he352;
aud[12355]=16'he33e;
aud[12356]=16'he32b;
aud[12357]=16'he318;
aud[12358]=16'he305;
aud[12359]=16'he2f2;
aud[12360]=16'he2df;
aud[12361]=16'he2cc;
aud[12362]=16'he2b9;
aud[12363]=16'he2a5;
aud[12364]=16'he292;
aud[12365]=16'he27f;
aud[12366]=16'he26c;
aud[12367]=16'he259;
aud[12368]=16'he246;
aud[12369]=16'he233;
aud[12370]=16'he220;
aud[12371]=16'he20d;
aud[12372]=16'he1fa;
aud[12373]=16'he1e8;
aud[12374]=16'he1d5;
aud[12375]=16'he1c2;
aud[12376]=16'he1af;
aud[12377]=16'he19c;
aud[12378]=16'he189;
aud[12379]=16'he176;
aud[12380]=16'he163;
aud[12381]=16'he151;
aud[12382]=16'he13e;
aud[12383]=16'he12b;
aud[12384]=16'he118;
aud[12385]=16'he105;
aud[12386]=16'he0f3;
aud[12387]=16'he0e0;
aud[12388]=16'he0cd;
aud[12389]=16'he0ba;
aud[12390]=16'he0a8;
aud[12391]=16'he095;
aud[12392]=16'he082;
aud[12393]=16'he070;
aud[12394]=16'he05d;
aud[12395]=16'he04a;
aud[12396]=16'he038;
aud[12397]=16'he025;
aud[12398]=16'he013;
aud[12399]=16'he000;
aud[12400]=16'hdfed;
aud[12401]=16'hdfdb;
aud[12402]=16'hdfc8;
aud[12403]=16'hdfb6;
aud[12404]=16'hdfa3;
aud[12405]=16'hdf91;
aud[12406]=16'hdf7e;
aud[12407]=16'hdf6c;
aud[12408]=16'hdf59;
aud[12409]=16'hdf47;
aud[12410]=16'hdf35;
aud[12411]=16'hdf22;
aud[12412]=16'hdf10;
aud[12413]=16'hdefd;
aud[12414]=16'hdeeb;
aud[12415]=16'hded9;
aud[12416]=16'hdec6;
aud[12417]=16'hdeb4;
aud[12418]=16'hdea2;
aud[12419]=16'hde8f;
aud[12420]=16'hde7d;
aud[12421]=16'hde6b;
aud[12422]=16'hde59;
aud[12423]=16'hde46;
aud[12424]=16'hde34;
aud[12425]=16'hde22;
aud[12426]=16'hde10;
aud[12427]=16'hddfe;
aud[12428]=16'hddeb;
aud[12429]=16'hddd9;
aud[12430]=16'hddc7;
aud[12431]=16'hddb5;
aud[12432]=16'hdda3;
aud[12433]=16'hdd91;
aud[12434]=16'hdd7f;
aud[12435]=16'hdd6d;
aud[12436]=16'hdd5b;
aud[12437]=16'hdd49;
aud[12438]=16'hdd37;
aud[12439]=16'hdd25;
aud[12440]=16'hdd13;
aud[12441]=16'hdd01;
aud[12442]=16'hdcef;
aud[12443]=16'hdcdd;
aud[12444]=16'hdccb;
aud[12445]=16'hdcb9;
aud[12446]=16'hdca7;
aud[12447]=16'hdc95;
aud[12448]=16'hdc83;
aud[12449]=16'hdc72;
aud[12450]=16'hdc60;
aud[12451]=16'hdc4e;
aud[12452]=16'hdc3c;
aud[12453]=16'hdc2a;
aud[12454]=16'hdc19;
aud[12455]=16'hdc07;
aud[12456]=16'hdbf5;
aud[12457]=16'hdbe3;
aud[12458]=16'hdbd2;
aud[12459]=16'hdbc0;
aud[12460]=16'hdbae;
aud[12461]=16'hdb9d;
aud[12462]=16'hdb8b;
aud[12463]=16'hdb79;
aud[12464]=16'hdb68;
aud[12465]=16'hdb56;
aud[12466]=16'hdb45;
aud[12467]=16'hdb33;
aud[12468]=16'hdb22;
aud[12469]=16'hdb10;
aud[12470]=16'hdaff;
aud[12471]=16'hdaed;
aud[12472]=16'hdadc;
aud[12473]=16'hdaca;
aud[12474]=16'hdab9;
aud[12475]=16'hdaa7;
aud[12476]=16'hda96;
aud[12477]=16'hda84;
aud[12478]=16'hda73;
aud[12479]=16'hda62;
aud[12480]=16'hda50;
aud[12481]=16'hda3f;
aud[12482]=16'hda2e;
aud[12483]=16'hda1c;
aud[12484]=16'hda0b;
aud[12485]=16'hd9fa;
aud[12486]=16'hd9e9;
aud[12487]=16'hd9d7;
aud[12488]=16'hd9c6;
aud[12489]=16'hd9b5;
aud[12490]=16'hd9a4;
aud[12491]=16'hd993;
aud[12492]=16'hd982;
aud[12493]=16'hd970;
aud[12494]=16'hd95f;
aud[12495]=16'hd94e;
aud[12496]=16'hd93d;
aud[12497]=16'hd92c;
aud[12498]=16'hd91b;
aud[12499]=16'hd90a;
aud[12500]=16'hd8f9;
aud[12501]=16'hd8e8;
aud[12502]=16'hd8d7;
aud[12503]=16'hd8c6;
aud[12504]=16'hd8b5;
aud[12505]=16'hd8a4;
aud[12506]=16'hd893;
aud[12507]=16'hd882;
aud[12508]=16'hd872;
aud[12509]=16'hd861;
aud[12510]=16'hd850;
aud[12511]=16'hd83f;
aud[12512]=16'hd82e;
aud[12513]=16'hd81e;
aud[12514]=16'hd80d;
aud[12515]=16'hd7fc;
aud[12516]=16'hd7eb;
aud[12517]=16'hd7db;
aud[12518]=16'hd7ca;
aud[12519]=16'hd7b9;
aud[12520]=16'hd7a9;
aud[12521]=16'hd798;
aud[12522]=16'hd787;
aud[12523]=16'hd777;
aud[12524]=16'hd766;
aud[12525]=16'hd756;
aud[12526]=16'hd745;
aud[12527]=16'hd734;
aud[12528]=16'hd724;
aud[12529]=16'hd713;
aud[12530]=16'hd703;
aud[12531]=16'hd6f2;
aud[12532]=16'hd6e2;
aud[12533]=16'hd6d2;
aud[12534]=16'hd6c1;
aud[12535]=16'hd6b1;
aud[12536]=16'hd6a0;
aud[12537]=16'hd690;
aud[12538]=16'hd680;
aud[12539]=16'hd66f;
aud[12540]=16'hd65f;
aud[12541]=16'hd64f;
aud[12542]=16'hd63f;
aud[12543]=16'hd62e;
aud[12544]=16'hd61e;
aud[12545]=16'hd60e;
aud[12546]=16'hd5fe;
aud[12547]=16'hd5ee;
aud[12548]=16'hd5dd;
aud[12549]=16'hd5cd;
aud[12550]=16'hd5bd;
aud[12551]=16'hd5ad;
aud[12552]=16'hd59d;
aud[12553]=16'hd58d;
aud[12554]=16'hd57d;
aud[12555]=16'hd56d;
aud[12556]=16'hd55d;
aud[12557]=16'hd54d;
aud[12558]=16'hd53d;
aud[12559]=16'hd52d;
aud[12560]=16'hd51d;
aud[12561]=16'hd50d;
aud[12562]=16'hd4fd;
aud[12563]=16'hd4ed;
aud[12564]=16'hd4de;
aud[12565]=16'hd4ce;
aud[12566]=16'hd4be;
aud[12567]=16'hd4ae;
aud[12568]=16'hd49e;
aud[12569]=16'hd48f;
aud[12570]=16'hd47f;
aud[12571]=16'hd46f;
aud[12572]=16'hd45f;
aud[12573]=16'hd450;
aud[12574]=16'hd440;
aud[12575]=16'hd430;
aud[12576]=16'hd421;
aud[12577]=16'hd411;
aud[12578]=16'hd402;
aud[12579]=16'hd3f2;
aud[12580]=16'hd3e2;
aud[12581]=16'hd3d3;
aud[12582]=16'hd3c3;
aud[12583]=16'hd3b4;
aud[12584]=16'hd3a4;
aud[12585]=16'hd395;
aud[12586]=16'hd386;
aud[12587]=16'hd376;
aud[12588]=16'hd367;
aud[12589]=16'hd357;
aud[12590]=16'hd348;
aud[12591]=16'hd339;
aud[12592]=16'hd329;
aud[12593]=16'hd31a;
aud[12594]=16'hd30b;
aud[12595]=16'hd2fc;
aud[12596]=16'hd2ec;
aud[12597]=16'hd2dd;
aud[12598]=16'hd2ce;
aud[12599]=16'hd2bf;
aud[12600]=16'hd2b0;
aud[12601]=16'hd2a0;
aud[12602]=16'hd291;
aud[12603]=16'hd282;
aud[12604]=16'hd273;
aud[12605]=16'hd264;
aud[12606]=16'hd255;
aud[12607]=16'hd246;
aud[12608]=16'hd237;
aud[12609]=16'hd228;
aud[12610]=16'hd219;
aud[12611]=16'hd20a;
aud[12612]=16'hd1fb;
aud[12613]=16'hd1ec;
aud[12614]=16'hd1de;
aud[12615]=16'hd1cf;
aud[12616]=16'hd1c0;
aud[12617]=16'hd1b1;
aud[12618]=16'hd1a2;
aud[12619]=16'hd193;
aud[12620]=16'hd185;
aud[12621]=16'hd176;
aud[12622]=16'hd167;
aud[12623]=16'hd159;
aud[12624]=16'hd14a;
aud[12625]=16'hd13b;
aud[12626]=16'hd12d;
aud[12627]=16'hd11e;
aud[12628]=16'hd10f;
aud[12629]=16'hd101;
aud[12630]=16'hd0f2;
aud[12631]=16'hd0e4;
aud[12632]=16'hd0d5;
aud[12633]=16'hd0c7;
aud[12634]=16'hd0b8;
aud[12635]=16'hd0aa;
aud[12636]=16'hd09b;
aud[12637]=16'hd08d;
aud[12638]=16'hd07f;
aud[12639]=16'hd070;
aud[12640]=16'hd062;
aud[12641]=16'hd054;
aud[12642]=16'hd045;
aud[12643]=16'hd037;
aud[12644]=16'hd029;
aud[12645]=16'hd01b;
aud[12646]=16'hd00c;
aud[12647]=16'hcffe;
aud[12648]=16'hcff0;
aud[12649]=16'hcfe2;
aud[12650]=16'hcfd4;
aud[12651]=16'hcfc6;
aud[12652]=16'hcfb8;
aud[12653]=16'hcfa9;
aud[12654]=16'hcf9b;
aud[12655]=16'hcf8d;
aud[12656]=16'hcf7f;
aud[12657]=16'hcf71;
aud[12658]=16'hcf63;
aud[12659]=16'hcf56;
aud[12660]=16'hcf48;
aud[12661]=16'hcf3a;
aud[12662]=16'hcf2c;
aud[12663]=16'hcf1e;
aud[12664]=16'hcf10;
aud[12665]=16'hcf02;
aud[12666]=16'hcef5;
aud[12667]=16'hcee7;
aud[12668]=16'hced9;
aud[12669]=16'hcecb;
aud[12670]=16'hcebe;
aud[12671]=16'hceb0;
aud[12672]=16'hcea2;
aud[12673]=16'hce95;
aud[12674]=16'hce87;
aud[12675]=16'hce79;
aud[12676]=16'hce6c;
aud[12677]=16'hce5e;
aud[12678]=16'hce51;
aud[12679]=16'hce43;
aud[12680]=16'hce36;
aud[12681]=16'hce28;
aud[12682]=16'hce1b;
aud[12683]=16'hce0d;
aud[12684]=16'hce00;
aud[12685]=16'hcdf3;
aud[12686]=16'hcde5;
aud[12687]=16'hcdd8;
aud[12688]=16'hcdcb;
aud[12689]=16'hcdbd;
aud[12690]=16'hcdb0;
aud[12691]=16'hcda3;
aud[12692]=16'hcd96;
aud[12693]=16'hcd88;
aud[12694]=16'hcd7b;
aud[12695]=16'hcd6e;
aud[12696]=16'hcd61;
aud[12697]=16'hcd54;
aud[12698]=16'hcd47;
aud[12699]=16'hcd3a;
aud[12700]=16'hcd2d;
aud[12701]=16'hcd20;
aud[12702]=16'hcd13;
aud[12703]=16'hcd06;
aud[12704]=16'hccf9;
aud[12705]=16'hccec;
aud[12706]=16'hccdf;
aud[12707]=16'hccd2;
aud[12708]=16'hccc5;
aud[12709]=16'hccb8;
aud[12710]=16'hccab;
aud[12711]=16'hcc9f;
aud[12712]=16'hcc92;
aud[12713]=16'hcc85;
aud[12714]=16'hcc78;
aud[12715]=16'hcc6c;
aud[12716]=16'hcc5f;
aud[12717]=16'hcc52;
aud[12718]=16'hcc46;
aud[12719]=16'hcc39;
aud[12720]=16'hcc2c;
aud[12721]=16'hcc20;
aud[12722]=16'hcc13;
aud[12723]=16'hcc07;
aud[12724]=16'hcbfa;
aud[12725]=16'hcbee;
aud[12726]=16'hcbe1;
aud[12727]=16'hcbd5;
aud[12728]=16'hcbc9;
aud[12729]=16'hcbbc;
aud[12730]=16'hcbb0;
aud[12731]=16'hcba3;
aud[12732]=16'hcb97;
aud[12733]=16'hcb8b;
aud[12734]=16'hcb7f;
aud[12735]=16'hcb72;
aud[12736]=16'hcb66;
aud[12737]=16'hcb5a;
aud[12738]=16'hcb4e;
aud[12739]=16'hcb42;
aud[12740]=16'hcb35;
aud[12741]=16'hcb29;
aud[12742]=16'hcb1d;
aud[12743]=16'hcb11;
aud[12744]=16'hcb05;
aud[12745]=16'hcaf9;
aud[12746]=16'hcaed;
aud[12747]=16'hcae1;
aud[12748]=16'hcad5;
aud[12749]=16'hcac9;
aud[12750]=16'hcabd;
aud[12751]=16'hcab1;
aud[12752]=16'hcaa6;
aud[12753]=16'hca9a;
aud[12754]=16'hca8e;
aud[12755]=16'hca82;
aud[12756]=16'hca76;
aud[12757]=16'hca6b;
aud[12758]=16'hca5f;
aud[12759]=16'hca53;
aud[12760]=16'hca48;
aud[12761]=16'hca3c;
aud[12762]=16'hca30;
aud[12763]=16'hca25;
aud[12764]=16'hca19;
aud[12765]=16'hca0e;
aud[12766]=16'hca02;
aud[12767]=16'hc9f7;
aud[12768]=16'hc9eb;
aud[12769]=16'hc9e0;
aud[12770]=16'hc9d4;
aud[12771]=16'hc9c9;
aud[12772]=16'hc9bd;
aud[12773]=16'hc9b2;
aud[12774]=16'hc9a7;
aud[12775]=16'hc99b;
aud[12776]=16'hc990;
aud[12777]=16'hc985;
aud[12778]=16'hc97a;
aud[12779]=16'hc96e;
aud[12780]=16'hc963;
aud[12781]=16'hc958;
aud[12782]=16'hc94d;
aud[12783]=16'hc942;
aud[12784]=16'hc937;
aud[12785]=16'hc92c;
aud[12786]=16'hc920;
aud[12787]=16'hc915;
aud[12788]=16'hc90a;
aud[12789]=16'hc8ff;
aud[12790]=16'hc8f5;
aud[12791]=16'hc8ea;
aud[12792]=16'hc8df;
aud[12793]=16'hc8d4;
aud[12794]=16'hc8c9;
aud[12795]=16'hc8be;
aud[12796]=16'hc8b3;
aud[12797]=16'hc8a9;
aud[12798]=16'hc89e;
aud[12799]=16'hc893;
aud[12800]=16'hc888;
aud[12801]=16'hc87e;
aud[12802]=16'hc873;
aud[12803]=16'hc868;
aud[12804]=16'hc85e;
aud[12805]=16'hc853;
aud[12806]=16'hc849;
aud[12807]=16'hc83e;
aud[12808]=16'hc834;
aud[12809]=16'hc829;
aud[12810]=16'hc81f;
aud[12811]=16'hc814;
aud[12812]=16'hc80a;
aud[12813]=16'hc7ff;
aud[12814]=16'hc7f5;
aud[12815]=16'hc7eb;
aud[12816]=16'hc7e0;
aud[12817]=16'hc7d6;
aud[12818]=16'hc7cc;
aud[12819]=16'hc7c1;
aud[12820]=16'hc7b7;
aud[12821]=16'hc7ad;
aud[12822]=16'hc7a3;
aud[12823]=16'hc799;
aud[12824]=16'hc78f;
aud[12825]=16'hc785;
aud[12826]=16'hc77a;
aud[12827]=16'hc770;
aud[12828]=16'hc766;
aud[12829]=16'hc75c;
aud[12830]=16'hc752;
aud[12831]=16'hc748;
aud[12832]=16'hc73f;
aud[12833]=16'hc735;
aud[12834]=16'hc72b;
aud[12835]=16'hc721;
aud[12836]=16'hc717;
aud[12837]=16'hc70d;
aud[12838]=16'hc703;
aud[12839]=16'hc6fa;
aud[12840]=16'hc6f0;
aud[12841]=16'hc6e6;
aud[12842]=16'hc6dd;
aud[12843]=16'hc6d3;
aud[12844]=16'hc6c9;
aud[12845]=16'hc6c0;
aud[12846]=16'hc6b6;
aud[12847]=16'hc6ad;
aud[12848]=16'hc6a3;
aud[12849]=16'hc69a;
aud[12850]=16'hc690;
aud[12851]=16'hc687;
aud[12852]=16'hc67d;
aud[12853]=16'hc674;
aud[12854]=16'hc66b;
aud[12855]=16'hc661;
aud[12856]=16'hc658;
aud[12857]=16'hc64f;
aud[12858]=16'hc645;
aud[12859]=16'hc63c;
aud[12860]=16'hc633;
aud[12861]=16'hc62a;
aud[12862]=16'hc620;
aud[12863]=16'hc617;
aud[12864]=16'hc60e;
aud[12865]=16'hc605;
aud[12866]=16'hc5fc;
aud[12867]=16'hc5f3;
aud[12868]=16'hc5ea;
aud[12869]=16'hc5e1;
aud[12870]=16'hc5d8;
aud[12871]=16'hc5cf;
aud[12872]=16'hc5c6;
aud[12873]=16'hc5bd;
aud[12874]=16'hc5b4;
aud[12875]=16'hc5ac;
aud[12876]=16'hc5a3;
aud[12877]=16'hc59a;
aud[12878]=16'hc591;
aud[12879]=16'hc588;
aud[12880]=16'hc580;
aud[12881]=16'hc577;
aud[12882]=16'hc56e;
aud[12883]=16'hc566;
aud[12884]=16'hc55d;
aud[12885]=16'hc555;
aud[12886]=16'hc54c;
aud[12887]=16'hc544;
aud[12888]=16'hc53b;
aud[12889]=16'hc533;
aud[12890]=16'hc52a;
aud[12891]=16'hc522;
aud[12892]=16'hc519;
aud[12893]=16'hc511;
aud[12894]=16'hc509;
aud[12895]=16'hc500;
aud[12896]=16'hc4f8;
aud[12897]=16'hc4f0;
aud[12898]=16'hc4e7;
aud[12899]=16'hc4df;
aud[12900]=16'hc4d7;
aud[12901]=16'hc4cf;
aud[12902]=16'hc4c7;
aud[12903]=16'hc4bf;
aud[12904]=16'hc4b6;
aud[12905]=16'hc4ae;
aud[12906]=16'hc4a6;
aud[12907]=16'hc49e;
aud[12908]=16'hc496;
aud[12909]=16'hc48e;
aud[12910]=16'hc486;
aud[12911]=16'hc47f;
aud[12912]=16'hc477;
aud[12913]=16'hc46f;
aud[12914]=16'hc467;
aud[12915]=16'hc45f;
aud[12916]=16'hc457;
aud[12917]=16'hc450;
aud[12918]=16'hc448;
aud[12919]=16'hc440;
aud[12920]=16'hc439;
aud[12921]=16'hc431;
aud[12922]=16'hc429;
aud[12923]=16'hc422;
aud[12924]=16'hc41a;
aud[12925]=16'hc413;
aud[12926]=16'hc40b;
aud[12927]=16'hc404;
aud[12928]=16'hc3fc;
aud[12929]=16'hc3f5;
aud[12930]=16'hc3ed;
aud[12931]=16'hc3e6;
aud[12932]=16'hc3df;
aud[12933]=16'hc3d7;
aud[12934]=16'hc3d0;
aud[12935]=16'hc3c9;
aud[12936]=16'hc3c1;
aud[12937]=16'hc3ba;
aud[12938]=16'hc3b3;
aud[12939]=16'hc3ac;
aud[12940]=16'hc3a5;
aud[12941]=16'hc39d;
aud[12942]=16'hc396;
aud[12943]=16'hc38f;
aud[12944]=16'hc388;
aud[12945]=16'hc381;
aud[12946]=16'hc37a;
aud[12947]=16'hc373;
aud[12948]=16'hc36c;
aud[12949]=16'hc365;
aud[12950]=16'hc35f;
aud[12951]=16'hc358;
aud[12952]=16'hc351;
aud[12953]=16'hc34a;
aud[12954]=16'hc343;
aud[12955]=16'hc33d;
aud[12956]=16'hc336;
aud[12957]=16'hc32f;
aud[12958]=16'hc329;
aud[12959]=16'hc322;
aud[12960]=16'hc31b;
aud[12961]=16'hc315;
aud[12962]=16'hc30e;
aud[12963]=16'hc308;
aud[12964]=16'hc301;
aud[12965]=16'hc2fb;
aud[12966]=16'hc2f4;
aud[12967]=16'hc2ee;
aud[12968]=16'hc2e7;
aud[12969]=16'hc2e1;
aud[12970]=16'hc2db;
aud[12971]=16'hc2d4;
aud[12972]=16'hc2ce;
aud[12973]=16'hc2c8;
aud[12974]=16'hc2c1;
aud[12975]=16'hc2bb;
aud[12976]=16'hc2b5;
aud[12977]=16'hc2af;
aud[12978]=16'hc2a9;
aud[12979]=16'hc2a3;
aud[12980]=16'hc29d;
aud[12981]=16'hc297;
aud[12982]=16'hc291;
aud[12983]=16'hc28b;
aud[12984]=16'hc285;
aud[12985]=16'hc27f;
aud[12986]=16'hc279;
aud[12987]=16'hc273;
aud[12988]=16'hc26d;
aud[12989]=16'hc267;
aud[12990]=16'hc261;
aud[12991]=16'hc25c;
aud[12992]=16'hc256;
aud[12993]=16'hc250;
aud[12994]=16'hc24a;
aud[12995]=16'hc245;
aud[12996]=16'hc23f;
aud[12997]=16'hc239;
aud[12998]=16'hc234;
aud[12999]=16'hc22e;
aud[13000]=16'hc229;
aud[13001]=16'hc223;
aud[13002]=16'hc21e;
aud[13003]=16'hc218;
aud[13004]=16'hc213;
aud[13005]=16'hc20d;
aud[13006]=16'hc208;
aud[13007]=16'hc203;
aud[13008]=16'hc1fd;
aud[13009]=16'hc1f8;
aud[13010]=16'hc1f3;
aud[13011]=16'hc1ee;
aud[13012]=16'hc1e8;
aud[13013]=16'hc1e3;
aud[13014]=16'hc1de;
aud[13015]=16'hc1d9;
aud[13016]=16'hc1d4;
aud[13017]=16'hc1cf;
aud[13018]=16'hc1ca;
aud[13019]=16'hc1c5;
aud[13020]=16'hc1c0;
aud[13021]=16'hc1bb;
aud[13022]=16'hc1b6;
aud[13023]=16'hc1b1;
aud[13024]=16'hc1ac;
aud[13025]=16'hc1a7;
aud[13026]=16'hc1a2;
aud[13027]=16'hc19e;
aud[13028]=16'hc199;
aud[13029]=16'hc194;
aud[13030]=16'hc18f;
aud[13031]=16'hc18b;
aud[13032]=16'hc186;
aud[13033]=16'hc181;
aud[13034]=16'hc17d;
aud[13035]=16'hc178;
aud[13036]=16'hc174;
aud[13037]=16'hc16f;
aud[13038]=16'hc16b;
aud[13039]=16'hc166;
aud[13040]=16'hc162;
aud[13041]=16'hc15d;
aud[13042]=16'hc159;
aud[13043]=16'hc154;
aud[13044]=16'hc150;
aud[13045]=16'hc14c;
aud[13046]=16'hc147;
aud[13047]=16'hc143;
aud[13048]=16'hc13f;
aud[13049]=16'hc13b;
aud[13050]=16'hc137;
aud[13051]=16'hc133;
aud[13052]=16'hc12e;
aud[13053]=16'hc12a;
aud[13054]=16'hc126;
aud[13055]=16'hc122;
aud[13056]=16'hc11e;
aud[13057]=16'hc11a;
aud[13058]=16'hc116;
aud[13059]=16'hc112;
aud[13060]=16'hc10e;
aud[13061]=16'hc10b;
aud[13062]=16'hc107;
aud[13063]=16'hc103;
aud[13064]=16'hc0ff;
aud[13065]=16'hc0fb;
aud[13066]=16'hc0f8;
aud[13067]=16'hc0f4;
aud[13068]=16'hc0f0;
aud[13069]=16'hc0ed;
aud[13070]=16'hc0e9;
aud[13071]=16'hc0e5;
aud[13072]=16'hc0e2;
aud[13073]=16'hc0de;
aud[13074]=16'hc0db;
aud[13075]=16'hc0d7;
aud[13076]=16'hc0d4;
aud[13077]=16'hc0d0;
aud[13078]=16'hc0cd;
aud[13079]=16'hc0ca;
aud[13080]=16'hc0c6;
aud[13081]=16'hc0c3;
aud[13082]=16'hc0c0;
aud[13083]=16'hc0bd;
aud[13084]=16'hc0b9;
aud[13085]=16'hc0b6;
aud[13086]=16'hc0b3;
aud[13087]=16'hc0b0;
aud[13088]=16'hc0ad;
aud[13089]=16'hc0aa;
aud[13090]=16'hc0a6;
aud[13091]=16'hc0a3;
aud[13092]=16'hc0a0;
aud[13093]=16'hc09d;
aud[13094]=16'hc09b;
aud[13095]=16'hc098;
aud[13096]=16'hc095;
aud[13097]=16'hc092;
aud[13098]=16'hc08f;
aud[13099]=16'hc08c;
aud[13100]=16'hc089;
aud[13101]=16'hc087;
aud[13102]=16'hc084;
aud[13103]=16'hc081;
aud[13104]=16'hc07f;
aud[13105]=16'hc07c;
aud[13106]=16'hc079;
aud[13107]=16'hc077;
aud[13108]=16'hc074;
aud[13109]=16'hc072;
aud[13110]=16'hc06f;
aud[13111]=16'hc06d;
aud[13112]=16'hc06a;
aud[13113]=16'hc068;
aud[13114]=16'hc065;
aud[13115]=16'hc063;
aud[13116]=16'hc061;
aud[13117]=16'hc05e;
aud[13118]=16'hc05c;
aud[13119]=16'hc05a;
aud[13120]=16'hc058;
aud[13121]=16'hc055;
aud[13122]=16'hc053;
aud[13123]=16'hc051;
aud[13124]=16'hc04f;
aud[13125]=16'hc04d;
aud[13126]=16'hc04b;
aud[13127]=16'hc049;
aud[13128]=16'hc047;
aud[13129]=16'hc045;
aud[13130]=16'hc043;
aud[13131]=16'hc041;
aud[13132]=16'hc03f;
aud[13133]=16'hc03d;
aud[13134]=16'hc03b;
aud[13135]=16'hc039;
aud[13136]=16'hc038;
aud[13137]=16'hc036;
aud[13138]=16'hc034;
aud[13139]=16'hc033;
aud[13140]=16'hc031;
aud[13141]=16'hc02f;
aud[13142]=16'hc02e;
aud[13143]=16'hc02c;
aud[13144]=16'hc02a;
aud[13145]=16'hc029;
aud[13146]=16'hc027;
aud[13147]=16'hc026;
aud[13148]=16'hc024;
aud[13149]=16'hc023;
aud[13150]=16'hc022;
aud[13151]=16'hc020;
aud[13152]=16'hc01f;
aud[13153]=16'hc01e;
aud[13154]=16'hc01c;
aud[13155]=16'hc01b;
aud[13156]=16'hc01a;
aud[13157]=16'hc019;
aud[13158]=16'hc018;
aud[13159]=16'hc016;
aud[13160]=16'hc015;
aud[13161]=16'hc014;
aud[13162]=16'hc013;
aud[13163]=16'hc012;
aud[13164]=16'hc011;
aud[13165]=16'hc010;
aud[13166]=16'hc00f;
aud[13167]=16'hc00e;
aud[13168]=16'hc00d;
aud[13169]=16'hc00d;
aud[13170]=16'hc00c;
aud[13171]=16'hc00b;
aud[13172]=16'hc00a;
aud[13173]=16'hc009;
aud[13174]=16'hc009;
aud[13175]=16'hc008;
aud[13176]=16'hc007;
aud[13177]=16'hc007;
aud[13178]=16'hc006;
aud[13179]=16'hc006;
aud[13180]=16'hc005;
aud[13181]=16'hc005;
aud[13182]=16'hc004;
aud[13183]=16'hc004;
aud[13184]=16'hc003;
aud[13185]=16'hc003;
aud[13186]=16'hc002;
aud[13187]=16'hc002;
aud[13188]=16'hc002;
aud[13189]=16'hc001;
aud[13190]=16'hc001;
aud[13191]=16'hc001;
aud[13192]=16'hc001;
aud[13193]=16'hc001;
aud[13194]=16'hc000;
aud[13195]=16'hc000;
aud[13196]=16'hc000;
aud[13197]=16'hc000;
aud[13198]=16'hc000;
aud[13199]=16'hc000;
aud[13200]=16'hc000;
aud[13201]=16'hc000;
aud[13202]=16'hc000;
aud[13203]=16'hc000;
aud[13204]=16'hc000;
aud[13205]=16'hc001;
aud[13206]=16'hc001;
aud[13207]=16'hc001;
aud[13208]=16'hc001;
aud[13209]=16'hc001;
aud[13210]=16'hc002;
aud[13211]=16'hc002;
aud[13212]=16'hc002;
aud[13213]=16'hc003;
aud[13214]=16'hc003;
aud[13215]=16'hc004;
aud[13216]=16'hc004;
aud[13217]=16'hc005;
aud[13218]=16'hc005;
aud[13219]=16'hc006;
aud[13220]=16'hc006;
aud[13221]=16'hc007;
aud[13222]=16'hc007;
aud[13223]=16'hc008;
aud[13224]=16'hc009;
aud[13225]=16'hc009;
aud[13226]=16'hc00a;
aud[13227]=16'hc00b;
aud[13228]=16'hc00c;
aud[13229]=16'hc00d;
aud[13230]=16'hc00d;
aud[13231]=16'hc00e;
aud[13232]=16'hc00f;
aud[13233]=16'hc010;
aud[13234]=16'hc011;
aud[13235]=16'hc012;
aud[13236]=16'hc013;
aud[13237]=16'hc014;
aud[13238]=16'hc015;
aud[13239]=16'hc016;
aud[13240]=16'hc018;
aud[13241]=16'hc019;
aud[13242]=16'hc01a;
aud[13243]=16'hc01b;
aud[13244]=16'hc01c;
aud[13245]=16'hc01e;
aud[13246]=16'hc01f;
aud[13247]=16'hc020;
aud[13248]=16'hc022;
aud[13249]=16'hc023;
aud[13250]=16'hc024;
aud[13251]=16'hc026;
aud[13252]=16'hc027;
aud[13253]=16'hc029;
aud[13254]=16'hc02a;
aud[13255]=16'hc02c;
aud[13256]=16'hc02e;
aud[13257]=16'hc02f;
aud[13258]=16'hc031;
aud[13259]=16'hc033;
aud[13260]=16'hc034;
aud[13261]=16'hc036;
aud[13262]=16'hc038;
aud[13263]=16'hc039;
aud[13264]=16'hc03b;
aud[13265]=16'hc03d;
aud[13266]=16'hc03f;
aud[13267]=16'hc041;
aud[13268]=16'hc043;
aud[13269]=16'hc045;
aud[13270]=16'hc047;
aud[13271]=16'hc049;
aud[13272]=16'hc04b;
aud[13273]=16'hc04d;
aud[13274]=16'hc04f;
aud[13275]=16'hc051;
aud[13276]=16'hc053;
aud[13277]=16'hc055;
aud[13278]=16'hc058;
aud[13279]=16'hc05a;
aud[13280]=16'hc05c;
aud[13281]=16'hc05e;
aud[13282]=16'hc061;
aud[13283]=16'hc063;
aud[13284]=16'hc065;
aud[13285]=16'hc068;
aud[13286]=16'hc06a;
aud[13287]=16'hc06d;
aud[13288]=16'hc06f;
aud[13289]=16'hc072;
aud[13290]=16'hc074;
aud[13291]=16'hc077;
aud[13292]=16'hc079;
aud[13293]=16'hc07c;
aud[13294]=16'hc07f;
aud[13295]=16'hc081;
aud[13296]=16'hc084;
aud[13297]=16'hc087;
aud[13298]=16'hc089;
aud[13299]=16'hc08c;
aud[13300]=16'hc08f;
aud[13301]=16'hc092;
aud[13302]=16'hc095;
aud[13303]=16'hc098;
aud[13304]=16'hc09b;
aud[13305]=16'hc09d;
aud[13306]=16'hc0a0;
aud[13307]=16'hc0a3;
aud[13308]=16'hc0a6;
aud[13309]=16'hc0aa;
aud[13310]=16'hc0ad;
aud[13311]=16'hc0b0;
aud[13312]=16'hc0b3;
aud[13313]=16'hc0b6;
aud[13314]=16'hc0b9;
aud[13315]=16'hc0bd;
aud[13316]=16'hc0c0;
aud[13317]=16'hc0c3;
aud[13318]=16'hc0c6;
aud[13319]=16'hc0ca;
aud[13320]=16'hc0cd;
aud[13321]=16'hc0d0;
aud[13322]=16'hc0d4;
aud[13323]=16'hc0d7;
aud[13324]=16'hc0db;
aud[13325]=16'hc0de;
aud[13326]=16'hc0e2;
aud[13327]=16'hc0e5;
aud[13328]=16'hc0e9;
aud[13329]=16'hc0ed;
aud[13330]=16'hc0f0;
aud[13331]=16'hc0f4;
aud[13332]=16'hc0f8;
aud[13333]=16'hc0fb;
aud[13334]=16'hc0ff;
aud[13335]=16'hc103;
aud[13336]=16'hc107;
aud[13337]=16'hc10b;
aud[13338]=16'hc10e;
aud[13339]=16'hc112;
aud[13340]=16'hc116;
aud[13341]=16'hc11a;
aud[13342]=16'hc11e;
aud[13343]=16'hc122;
aud[13344]=16'hc126;
aud[13345]=16'hc12a;
aud[13346]=16'hc12e;
aud[13347]=16'hc133;
aud[13348]=16'hc137;
aud[13349]=16'hc13b;
aud[13350]=16'hc13f;
aud[13351]=16'hc143;
aud[13352]=16'hc147;
aud[13353]=16'hc14c;
aud[13354]=16'hc150;
aud[13355]=16'hc154;
aud[13356]=16'hc159;
aud[13357]=16'hc15d;
aud[13358]=16'hc162;
aud[13359]=16'hc166;
aud[13360]=16'hc16b;
aud[13361]=16'hc16f;
aud[13362]=16'hc174;
aud[13363]=16'hc178;
aud[13364]=16'hc17d;
aud[13365]=16'hc181;
aud[13366]=16'hc186;
aud[13367]=16'hc18b;
aud[13368]=16'hc18f;
aud[13369]=16'hc194;
aud[13370]=16'hc199;
aud[13371]=16'hc19e;
aud[13372]=16'hc1a2;
aud[13373]=16'hc1a7;
aud[13374]=16'hc1ac;
aud[13375]=16'hc1b1;
aud[13376]=16'hc1b6;
aud[13377]=16'hc1bb;
aud[13378]=16'hc1c0;
aud[13379]=16'hc1c5;
aud[13380]=16'hc1ca;
aud[13381]=16'hc1cf;
aud[13382]=16'hc1d4;
aud[13383]=16'hc1d9;
aud[13384]=16'hc1de;
aud[13385]=16'hc1e3;
aud[13386]=16'hc1e8;
aud[13387]=16'hc1ee;
aud[13388]=16'hc1f3;
aud[13389]=16'hc1f8;
aud[13390]=16'hc1fd;
aud[13391]=16'hc203;
aud[13392]=16'hc208;
aud[13393]=16'hc20d;
aud[13394]=16'hc213;
aud[13395]=16'hc218;
aud[13396]=16'hc21e;
aud[13397]=16'hc223;
aud[13398]=16'hc229;
aud[13399]=16'hc22e;
aud[13400]=16'hc234;
aud[13401]=16'hc239;
aud[13402]=16'hc23f;
aud[13403]=16'hc245;
aud[13404]=16'hc24a;
aud[13405]=16'hc250;
aud[13406]=16'hc256;
aud[13407]=16'hc25c;
aud[13408]=16'hc261;
aud[13409]=16'hc267;
aud[13410]=16'hc26d;
aud[13411]=16'hc273;
aud[13412]=16'hc279;
aud[13413]=16'hc27f;
aud[13414]=16'hc285;
aud[13415]=16'hc28b;
aud[13416]=16'hc291;
aud[13417]=16'hc297;
aud[13418]=16'hc29d;
aud[13419]=16'hc2a3;
aud[13420]=16'hc2a9;
aud[13421]=16'hc2af;
aud[13422]=16'hc2b5;
aud[13423]=16'hc2bb;
aud[13424]=16'hc2c1;
aud[13425]=16'hc2c8;
aud[13426]=16'hc2ce;
aud[13427]=16'hc2d4;
aud[13428]=16'hc2db;
aud[13429]=16'hc2e1;
aud[13430]=16'hc2e7;
aud[13431]=16'hc2ee;
aud[13432]=16'hc2f4;
aud[13433]=16'hc2fb;
aud[13434]=16'hc301;
aud[13435]=16'hc308;
aud[13436]=16'hc30e;
aud[13437]=16'hc315;
aud[13438]=16'hc31b;
aud[13439]=16'hc322;
aud[13440]=16'hc329;
aud[13441]=16'hc32f;
aud[13442]=16'hc336;
aud[13443]=16'hc33d;
aud[13444]=16'hc343;
aud[13445]=16'hc34a;
aud[13446]=16'hc351;
aud[13447]=16'hc358;
aud[13448]=16'hc35f;
aud[13449]=16'hc365;
aud[13450]=16'hc36c;
aud[13451]=16'hc373;
aud[13452]=16'hc37a;
aud[13453]=16'hc381;
aud[13454]=16'hc388;
aud[13455]=16'hc38f;
aud[13456]=16'hc396;
aud[13457]=16'hc39d;
aud[13458]=16'hc3a5;
aud[13459]=16'hc3ac;
aud[13460]=16'hc3b3;
aud[13461]=16'hc3ba;
aud[13462]=16'hc3c1;
aud[13463]=16'hc3c9;
aud[13464]=16'hc3d0;
aud[13465]=16'hc3d7;
aud[13466]=16'hc3df;
aud[13467]=16'hc3e6;
aud[13468]=16'hc3ed;
aud[13469]=16'hc3f5;
aud[13470]=16'hc3fc;
aud[13471]=16'hc404;
aud[13472]=16'hc40b;
aud[13473]=16'hc413;
aud[13474]=16'hc41a;
aud[13475]=16'hc422;
aud[13476]=16'hc429;
aud[13477]=16'hc431;
aud[13478]=16'hc439;
aud[13479]=16'hc440;
aud[13480]=16'hc448;
aud[13481]=16'hc450;
aud[13482]=16'hc457;
aud[13483]=16'hc45f;
aud[13484]=16'hc467;
aud[13485]=16'hc46f;
aud[13486]=16'hc477;
aud[13487]=16'hc47f;
aud[13488]=16'hc486;
aud[13489]=16'hc48e;
aud[13490]=16'hc496;
aud[13491]=16'hc49e;
aud[13492]=16'hc4a6;
aud[13493]=16'hc4ae;
aud[13494]=16'hc4b6;
aud[13495]=16'hc4bf;
aud[13496]=16'hc4c7;
aud[13497]=16'hc4cf;
aud[13498]=16'hc4d7;
aud[13499]=16'hc4df;
aud[13500]=16'hc4e7;
aud[13501]=16'hc4f0;
aud[13502]=16'hc4f8;
aud[13503]=16'hc500;
aud[13504]=16'hc509;
aud[13505]=16'hc511;
aud[13506]=16'hc519;
aud[13507]=16'hc522;
aud[13508]=16'hc52a;
aud[13509]=16'hc533;
aud[13510]=16'hc53b;
aud[13511]=16'hc544;
aud[13512]=16'hc54c;
aud[13513]=16'hc555;
aud[13514]=16'hc55d;
aud[13515]=16'hc566;
aud[13516]=16'hc56e;
aud[13517]=16'hc577;
aud[13518]=16'hc580;
aud[13519]=16'hc588;
aud[13520]=16'hc591;
aud[13521]=16'hc59a;
aud[13522]=16'hc5a3;
aud[13523]=16'hc5ac;
aud[13524]=16'hc5b4;
aud[13525]=16'hc5bd;
aud[13526]=16'hc5c6;
aud[13527]=16'hc5cf;
aud[13528]=16'hc5d8;
aud[13529]=16'hc5e1;
aud[13530]=16'hc5ea;
aud[13531]=16'hc5f3;
aud[13532]=16'hc5fc;
aud[13533]=16'hc605;
aud[13534]=16'hc60e;
aud[13535]=16'hc617;
aud[13536]=16'hc620;
aud[13537]=16'hc62a;
aud[13538]=16'hc633;
aud[13539]=16'hc63c;
aud[13540]=16'hc645;
aud[13541]=16'hc64f;
aud[13542]=16'hc658;
aud[13543]=16'hc661;
aud[13544]=16'hc66b;
aud[13545]=16'hc674;
aud[13546]=16'hc67d;
aud[13547]=16'hc687;
aud[13548]=16'hc690;
aud[13549]=16'hc69a;
aud[13550]=16'hc6a3;
aud[13551]=16'hc6ad;
aud[13552]=16'hc6b6;
aud[13553]=16'hc6c0;
aud[13554]=16'hc6c9;
aud[13555]=16'hc6d3;
aud[13556]=16'hc6dd;
aud[13557]=16'hc6e6;
aud[13558]=16'hc6f0;
aud[13559]=16'hc6fa;
aud[13560]=16'hc703;
aud[13561]=16'hc70d;
aud[13562]=16'hc717;
aud[13563]=16'hc721;
aud[13564]=16'hc72b;
aud[13565]=16'hc735;
aud[13566]=16'hc73f;
aud[13567]=16'hc748;
aud[13568]=16'hc752;
aud[13569]=16'hc75c;
aud[13570]=16'hc766;
aud[13571]=16'hc770;
aud[13572]=16'hc77a;
aud[13573]=16'hc785;
aud[13574]=16'hc78f;
aud[13575]=16'hc799;
aud[13576]=16'hc7a3;
aud[13577]=16'hc7ad;
aud[13578]=16'hc7b7;
aud[13579]=16'hc7c1;
aud[13580]=16'hc7cc;
aud[13581]=16'hc7d6;
aud[13582]=16'hc7e0;
aud[13583]=16'hc7eb;
aud[13584]=16'hc7f5;
aud[13585]=16'hc7ff;
aud[13586]=16'hc80a;
aud[13587]=16'hc814;
aud[13588]=16'hc81f;
aud[13589]=16'hc829;
aud[13590]=16'hc834;
aud[13591]=16'hc83e;
aud[13592]=16'hc849;
aud[13593]=16'hc853;
aud[13594]=16'hc85e;
aud[13595]=16'hc868;
aud[13596]=16'hc873;
aud[13597]=16'hc87e;
aud[13598]=16'hc888;
aud[13599]=16'hc893;
aud[13600]=16'hc89e;
aud[13601]=16'hc8a9;
aud[13602]=16'hc8b3;
aud[13603]=16'hc8be;
aud[13604]=16'hc8c9;
aud[13605]=16'hc8d4;
aud[13606]=16'hc8df;
aud[13607]=16'hc8ea;
aud[13608]=16'hc8f5;
aud[13609]=16'hc8ff;
aud[13610]=16'hc90a;
aud[13611]=16'hc915;
aud[13612]=16'hc920;
aud[13613]=16'hc92c;
aud[13614]=16'hc937;
aud[13615]=16'hc942;
aud[13616]=16'hc94d;
aud[13617]=16'hc958;
aud[13618]=16'hc963;
aud[13619]=16'hc96e;
aud[13620]=16'hc97a;
aud[13621]=16'hc985;
aud[13622]=16'hc990;
aud[13623]=16'hc99b;
aud[13624]=16'hc9a7;
aud[13625]=16'hc9b2;
aud[13626]=16'hc9bd;
aud[13627]=16'hc9c9;
aud[13628]=16'hc9d4;
aud[13629]=16'hc9e0;
aud[13630]=16'hc9eb;
aud[13631]=16'hc9f7;
aud[13632]=16'hca02;
aud[13633]=16'hca0e;
aud[13634]=16'hca19;
aud[13635]=16'hca25;
aud[13636]=16'hca30;
aud[13637]=16'hca3c;
aud[13638]=16'hca48;
aud[13639]=16'hca53;
aud[13640]=16'hca5f;
aud[13641]=16'hca6b;
aud[13642]=16'hca76;
aud[13643]=16'hca82;
aud[13644]=16'hca8e;
aud[13645]=16'hca9a;
aud[13646]=16'hcaa6;
aud[13647]=16'hcab1;
aud[13648]=16'hcabd;
aud[13649]=16'hcac9;
aud[13650]=16'hcad5;
aud[13651]=16'hcae1;
aud[13652]=16'hcaed;
aud[13653]=16'hcaf9;
aud[13654]=16'hcb05;
aud[13655]=16'hcb11;
aud[13656]=16'hcb1d;
aud[13657]=16'hcb29;
aud[13658]=16'hcb35;
aud[13659]=16'hcb42;
aud[13660]=16'hcb4e;
aud[13661]=16'hcb5a;
aud[13662]=16'hcb66;
aud[13663]=16'hcb72;
aud[13664]=16'hcb7f;
aud[13665]=16'hcb8b;
aud[13666]=16'hcb97;
aud[13667]=16'hcba3;
aud[13668]=16'hcbb0;
aud[13669]=16'hcbbc;
aud[13670]=16'hcbc9;
aud[13671]=16'hcbd5;
aud[13672]=16'hcbe1;
aud[13673]=16'hcbee;
aud[13674]=16'hcbfa;
aud[13675]=16'hcc07;
aud[13676]=16'hcc13;
aud[13677]=16'hcc20;
aud[13678]=16'hcc2c;
aud[13679]=16'hcc39;
aud[13680]=16'hcc46;
aud[13681]=16'hcc52;
aud[13682]=16'hcc5f;
aud[13683]=16'hcc6c;
aud[13684]=16'hcc78;
aud[13685]=16'hcc85;
aud[13686]=16'hcc92;
aud[13687]=16'hcc9f;
aud[13688]=16'hccab;
aud[13689]=16'hccb8;
aud[13690]=16'hccc5;
aud[13691]=16'hccd2;
aud[13692]=16'hccdf;
aud[13693]=16'hccec;
aud[13694]=16'hccf9;
aud[13695]=16'hcd06;
aud[13696]=16'hcd13;
aud[13697]=16'hcd20;
aud[13698]=16'hcd2d;
aud[13699]=16'hcd3a;
aud[13700]=16'hcd47;
aud[13701]=16'hcd54;
aud[13702]=16'hcd61;
aud[13703]=16'hcd6e;
aud[13704]=16'hcd7b;
aud[13705]=16'hcd88;
aud[13706]=16'hcd96;
aud[13707]=16'hcda3;
aud[13708]=16'hcdb0;
aud[13709]=16'hcdbd;
aud[13710]=16'hcdcb;
aud[13711]=16'hcdd8;
aud[13712]=16'hcde5;
aud[13713]=16'hcdf3;
aud[13714]=16'hce00;
aud[13715]=16'hce0d;
aud[13716]=16'hce1b;
aud[13717]=16'hce28;
aud[13718]=16'hce36;
aud[13719]=16'hce43;
aud[13720]=16'hce51;
aud[13721]=16'hce5e;
aud[13722]=16'hce6c;
aud[13723]=16'hce79;
aud[13724]=16'hce87;
aud[13725]=16'hce95;
aud[13726]=16'hcea2;
aud[13727]=16'hceb0;
aud[13728]=16'hcebe;
aud[13729]=16'hcecb;
aud[13730]=16'hced9;
aud[13731]=16'hcee7;
aud[13732]=16'hcef5;
aud[13733]=16'hcf02;
aud[13734]=16'hcf10;
aud[13735]=16'hcf1e;
aud[13736]=16'hcf2c;
aud[13737]=16'hcf3a;
aud[13738]=16'hcf48;
aud[13739]=16'hcf56;
aud[13740]=16'hcf63;
aud[13741]=16'hcf71;
aud[13742]=16'hcf7f;
aud[13743]=16'hcf8d;
aud[13744]=16'hcf9b;
aud[13745]=16'hcfa9;
aud[13746]=16'hcfb8;
aud[13747]=16'hcfc6;
aud[13748]=16'hcfd4;
aud[13749]=16'hcfe2;
aud[13750]=16'hcff0;
aud[13751]=16'hcffe;
aud[13752]=16'hd00c;
aud[13753]=16'hd01b;
aud[13754]=16'hd029;
aud[13755]=16'hd037;
aud[13756]=16'hd045;
aud[13757]=16'hd054;
aud[13758]=16'hd062;
aud[13759]=16'hd070;
aud[13760]=16'hd07f;
aud[13761]=16'hd08d;
aud[13762]=16'hd09b;
aud[13763]=16'hd0aa;
aud[13764]=16'hd0b8;
aud[13765]=16'hd0c7;
aud[13766]=16'hd0d5;
aud[13767]=16'hd0e4;
aud[13768]=16'hd0f2;
aud[13769]=16'hd101;
aud[13770]=16'hd10f;
aud[13771]=16'hd11e;
aud[13772]=16'hd12d;
aud[13773]=16'hd13b;
aud[13774]=16'hd14a;
aud[13775]=16'hd159;
aud[13776]=16'hd167;
aud[13777]=16'hd176;
aud[13778]=16'hd185;
aud[13779]=16'hd193;
aud[13780]=16'hd1a2;
aud[13781]=16'hd1b1;
aud[13782]=16'hd1c0;
aud[13783]=16'hd1cf;
aud[13784]=16'hd1de;
aud[13785]=16'hd1ec;
aud[13786]=16'hd1fb;
aud[13787]=16'hd20a;
aud[13788]=16'hd219;
aud[13789]=16'hd228;
aud[13790]=16'hd237;
aud[13791]=16'hd246;
aud[13792]=16'hd255;
aud[13793]=16'hd264;
aud[13794]=16'hd273;
aud[13795]=16'hd282;
aud[13796]=16'hd291;
aud[13797]=16'hd2a0;
aud[13798]=16'hd2b0;
aud[13799]=16'hd2bf;
aud[13800]=16'hd2ce;
aud[13801]=16'hd2dd;
aud[13802]=16'hd2ec;
aud[13803]=16'hd2fc;
aud[13804]=16'hd30b;
aud[13805]=16'hd31a;
aud[13806]=16'hd329;
aud[13807]=16'hd339;
aud[13808]=16'hd348;
aud[13809]=16'hd357;
aud[13810]=16'hd367;
aud[13811]=16'hd376;
aud[13812]=16'hd386;
aud[13813]=16'hd395;
aud[13814]=16'hd3a4;
aud[13815]=16'hd3b4;
aud[13816]=16'hd3c3;
aud[13817]=16'hd3d3;
aud[13818]=16'hd3e2;
aud[13819]=16'hd3f2;
aud[13820]=16'hd402;
aud[13821]=16'hd411;
aud[13822]=16'hd421;
aud[13823]=16'hd430;
aud[13824]=16'hd440;
aud[13825]=16'hd450;
aud[13826]=16'hd45f;
aud[13827]=16'hd46f;
aud[13828]=16'hd47f;
aud[13829]=16'hd48f;
aud[13830]=16'hd49e;
aud[13831]=16'hd4ae;
aud[13832]=16'hd4be;
aud[13833]=16'hd4ce;
aud[13834]=16'hd4de;
aud[13835]=16'hd4ed;
aud[13836]=16'hd4fd;
aud[13837]=16'hd50d;
aud[13838]=16'hd51d;
aud[13839]=16'hd52d;
aud[13840]=16'hd53d;
aud[13841]=16'hd54d;
aud[13842]=16'hd55d;
aud[13843]=16'hd56d;
aud[13844]=16'hd57d;
aud[13845]=16'hd58d;
aud[13846]=16'hd59d;
aud[13847]=16'hd5ad;
aud[13848]=16'hd5bd;
aud[13849]=16'hd5cd;
aud[13850]=16'hd5dd;
aud[13851]=16'hd5ee;
aud[13852]=16'hd5fe;
aud[13853]=16'hd60e;
aud[13854]=16'hd61e;
aud[13855]=16'hd62e;
aud[13856]=16'hd63f;
aud[13857]=16'hd64f;
aud[13858]=16'hd65f;
aud[13859]=16'hd66f;
aud[13860]=16'hd680;
aud[13861]=16'hd690;
aud[13862]=16'hd6a0;
aud[13863]=16'hd6b1;
aud[13864]=16'hd6c1;
aud[13865]=16'hd6d2;
aud[13866]=16'hd6e2;
aud[13867]=16'hd6f2;
aud[13868]=16'hd703;
aud[13869]=16'hd713;
aud[13870]=16'hd724;
aud[13871]=16'hd734;
aud[13872]=16'hd745;
aud[13873]=16'hd756;
aud[13874]=16'hd766;
aud[13875]=16'hd777;
aud[13876]=16'hd787;
aud[13877]=16'hd798;
aud[13878]=16'hd7a9;
aud[13879]=16'hd7b9;
aud[13880]=16'hd7ca;
aud[13881]=16'hd7db;
aud[13882]=16'hd7eb;
aud[13883]=16'hd7fc;
aud[13884]=16'hd80d;
aud[13885]=16'hd81e;
aud[13886]=16'hd82e;
aud[13887]=16'hd83f;
aud[13888]=16'hd850;
aud[13889]=16'hd861;
aud[13890]=16'hd872;
aud[13891]=16'hd882;
aud[13892]=16'hd893;
aud[13893]=16'hd8a4;
aud[13894]=16'hd8b5;
aud[13895]=16'hd8c6;
aud[13896]=16'hd8d7;
aud[13897]=16'hd8e8;
aud[13898]=16'hd8f9;
aud[13899]=16'hd90a;
aud[13900]=16'hd91b;
aud[13901]=16'hd92c;
aud[13902]=16'hd93d;
aud[13903]=16'hd94e;
aud[13904]=16'hd95f;
aud[13905]=16'hd970;
aud[13906]=16'hd982;
aud[13907]=16'hd993;
aud[13908]=16'hd9a4;
aud[13909]=16'hd9b5;
aud[13910]=16'hd9c6;
aud[13911]=16'hd9d7;
aud[13912]=16'hd9e9;
aud[13913]=16'hd9fa;
aud[13914]=16'hda0b;
aud[13915]=16'hda1c;
aud[13916]=16'hda2e;
aud[13917]=16'hda3f;
aud[13918]=16'hda50;
aud[13919]=16'hda62;
aud[13920]=16'hda73;
aud[13921]=16'hda84;
aud[13922]=16'hda96;
aud[13923]=16'hdaa7;
aud[13924]=16'hdab9;
aud[13925]=16'hdaca;
aud[13926]=16'hdadc;
aud[13927]=16'hdaed;
aud[13928]=16'hdaff;
aud[13929]=16'hdb10;
aud[13930]=16'hdb22;
aud[13931]=16'hdb33;
aud[13932]=16'hdb45;
aud[13933]=16'hdb56;
aud[13934]=16'hdb68;
aud[13935]=16'hdb79;
aud[13936]=16'hdb8b;
aud[13937]=16'hdb9d;
aud[13938]=16'hdbae;
aud[13939]=16'hdbc0;
aud[13940]=16'hdbd2;
aud[13941]=16'hdbe3;
aud[13942]=16'hdbf5;
aud[13943]=16'hdc07;
aud[13944]=16'hdc19;
aud[13945]=16'hdc2a;
aud[13946]=16'hdc3c;
aud[13947]=16'hdc4e;
aud[13948]=16'hdc60;
aud[13949]=16'hdc72;
aud[13950]=16'hdc83;
aud[13951]=16'hdc95;
aud[13952]=16'hdca7;
aud[13953]=16'hdcb9;
aud[13954]=16'hdccb;
aud[13955]=16'hdcdd;
aud[13956]=16'hdcef;
aud[13957]=16'hdd01;
aud[13958]=16'hdd13;
aud[13959]=16'hdd25;
aud[13960]=16'hdd37;
aud[13961]=16'hdd49;
aud[13962]=16'hdd5b;
aud[13963]=16'hdd6d;
aud[13964]=16'hdd7f;
aud[13965]=16'hdd91;
aud[13966]=16'hdda3;
aud[13967]=16'hddb5;
aud[13968]=16'hddc7;
aud[13969]=16'hddd9;
aud[13970]=16'hddeb;
aud[13971]=16'hddfe;
aud[13972]=16'hde10;
aud[13973]=16'hde22;
aud[13974]=16'hde34;
aud[13975]=16'hde46;
aud[13976]=16'hde59;
aud[13977]=16'hde6b;
aud[13978]=16'hde7d;
aud[13979]=16'hde8f;
aud[13980]=16'hdea2;
aud[13981]=16'hdeb4;
aud[13982]=16'hdec6;
aud[13983]=16'hded9;
aud[13984]=16'hdeeb;
aud[13985]=16'hdefd;
aud[13986]=16'hdf10;
aud[13987]=16'hdf22;
aud[13988]=16'hdf35;
aud[13989]=16'hdf47;
aud[13990]=16'hdf59;
aud[13991]=16'hdf6c;
aud[13992]=16'hdf7e;
aud[13993]=16'hdf91;
aud[13994]=16'hdfa3;
aud[13995]=16'hdfb6;
aud[13996]=16'hdfc8;
aud[13997]=16'hdfdb;
aud[13998]=16'hdfed;
aud[13999]=16'he000;
aud[14000]=16'he013;
aud[14001]=16'he025;
aud[14002]=16'he038;
aud[14003]=16'he04a;
aud[14004]=16'he05d;
aud[14005]=16'he070;
aud[14006]=16'he082;
aud[14007]=16'he095;
aud[14008]=16'he0a8;
aud[14009]=16'he0ba;
aud[14010]=16'he0cd;
aud[14011]=16'he0e0;
aud[14012]=16'he0f3;
aud[14013]=16'he105;
aud[14014]=16'he118;
aud[14015]=16'he12b;
aud[14016]=16'he13e;
aud[14017]=16'he151;
aud[14018]=16'he163;
aud[14019]=16'he176;
aud[14020]=16'he189;
aud[14021]=16'he19c;
aud[14022]=16'he1af;
aud[14023]=16'he1c2;
aud[14024]=16'he1d5;
aud[14025]=16'he1e8;
aud[14026]=16'he1fa;
aud[14027]=16'he20d;
aud[14028]=16'he220;
aud[14029]=16'he233;
aud[14030]=16'he246;
aud[14031]=16'he259;
aud[14032]=16'he26c;
aud[14033]=16'he27f;
aud[14034]=16'he292;
aud[14035]=16'he2a5;
aud[14036]=16'he2b9;
aud[14037]=16'he2cc;
aud[14038]=16'he2df;
aud[14039]=16'he2f2;
aud[14040]=16'he305;
aud[14041]=16'he318;
aud[14042]=16'he32b;
aud[14043]=16'he33e;
aud[14044]=16'he352;
aud[14045]=16'he365;
aud[14046]=16'he378;
aud[14047]=16'he38b;
aud[14048]=16'he39e;
aud[14049]=16'he3b2;
aud[14050]=16'he3c5;
aud[14051]=16'he3d8;
aud[14052]=16'he3eb;
aud[14053]=16'he3ff;
aud[14054]=16'he412;
aud[14055]=16'he425;
aud[14056]=16'he438;
aud[14057]=16'he44c;
aud[14058]=16'he45f;
aud[14059]=16'he473;
aud[14060]=16'he486;
aud[14061]=16'he499;
aud[14062]=16'he4ad;
aud[14063]=16'he4c0;
aud[14064]=16'he4d3;
aud[14065]=16'he4e7;
aud[14066]=16'he4fa;
aud[14067]=16'he50e;
aud[14068]=16'he521;
aud[14069]=16'he535;
aud[14070]=16'he548;
aud[14071]=16'he55c;
aud[14072]=16'he56f;
aud[14073]=16'he583;
aud[14074]=16'he596;
aud[14075]=16'he5aa;
aud[14076]=16'he5bd;
aud[14077]=16'he5d1;
aud[14078]=16'he5e4;
aud[14079]=16'he5f8;
aud[14080]=16'he60c;
aud[14081]=16'he61f;
aud[14082]=16'he633;
aud[14083]=16'he646;
aud[14084]=16'he65a;
aud[14085]=16'he66e;
aud[14086]=16'he681;
aud[14087]=16'he695;
aud[14088]=16'he6a9;
aud[14089]=16'he6bd;
aud[14090]=16'he6d0;
aud[14091]=16'he6e4;
aud[14092]=16'he6f8;
aud[14093]=16'he70b;
aud[14094]=16'he71f;
aud[14095]=16'he733;
aud[14096]=16'he747;
aud[14097]=16'he75b;
aud[14098]=16'he76e;
aud[14099]=16'he782;
aud[14100]=16'he796;
aud[14101]=16'he7aa;
aud[14102]=16'he7be;
aud[14103]=16'he7d1;
aud[14104]=16'he7e5;
aud[14105]=16'he7f9;
aud[14106]=16'he80d;
aud[14107]=16'he821;
aud[14108]=16'he835;
aud[14109]=16'he849;
aud[14110]=16'he85d;
aud[14111]=16'he871;
aud[14112]=16'he885;
aud[14113]=16'he899;
aud[14114]=16'he8ad;
aud[14115]=16'he8c0;
aud[14116]=16'he8d4;
aud[14117]=16'he8e8;
aud[14118]=16'he8fc;
aud[14119]=16'he910;
aud[14120]=16'he925;
aud[14121]=16'he939;
aud[14122]=16'he94d;
aud[14123]=16'he961;
aud[14124]=16'he975;
aud[14125]=16'he989;
aud[14126]=16'he99d;
aud[14127]=16'he9b1;
aud[14128]=16'he9c5;
aud[14129]=16'he9d9;
aud[14130]=16'he9ed;
aud[14131]=16'hea01;
aud[14132]=16'hea16;
aud[14133]=16'hea2a;
aud[14134]=16'hea3e;
aud[14135]=16'hea52;
aud[14136]=16'hea66;
aud[14137]=16'hea7a;
aud[14138]=16'hea8f;
aud[14139]=16'heaa3;
aud[14140]=16'heab7;
aud[14141]=16'heacb;
aud[14142]=16'heae0;
aud[14143]=16'heaf4;
aud[14144]=16'heb08;
aud[14145]=16'heb1c;
aud[14146]=16'heb31;
aud[14147]=16'heb45;
aud[14148]=16'heb59;
aud[14149]=16'heb6e;
aud[14150]=16'heb82;
aud[14151]=16'heb96;
aud[14152]=16'hebab;
aud[14153]=16'hebbf;
aud[14154]=16'hebd3;
aud[14155]=16'hebe8;
aud[14156]=16'hebfc;
aud[14157]=16'hec10;
aud[14158]=16'hec25;
aud[14159]=16'hec39;
aud[14160]=16'hec4d;
aud[14161]=16'hec62;
aud[14162]=16'hec76;
aud[14163]=16'hec8b;
aud[14164]=16'hec9f;
aud[14165]=16'hecb4;
aud[14166]=16'hecc8;
aud[14167]=16'hecdd;
aud[14168]=16'hecf1;
aud[14169]=16'hed05;
aud[14170]=16'hed1a;
aud[14171]=16'hed2e;
aud[14172]=16'hed43;
aud[14173]=16'hed57;
aud[14174]=16'hed6c;
aud[14175]=16'hed81;
aud[14176]=16'hed95;
aud[14177]=16'hedaa;
aud[14178]=16'hedbe;
aud[14179]=16'hedd3;
aud[14180]=16'hede7;
aud[14181]=16'hedfc;
aud[14182]=16'hee10;
aud[14183]=16'hee25;
aud[14184]=16'hee3a;
aud[14185]=16'hee4e;
aud[14186]=16'hee63;
aud[14187]=16'hee77;
aud[14188]=16'hee8c;
aud[14189]=16'heea1;
aud[14190]=16'heeb5;
aud[14191]=16'heeca;
aud[14192]=16'heedf;
aud[14193]=16'heef3;
aud[14194]=16'hef08;
aud[14195]=16'hef1d;
aud[14196]=16'hef31;
aud[14197]=16'hef46;
aud[14198]=16'hef5b;
aud[14199]=16'hef70;
aud[14200]=16'hef84;
aud[14201]=16'hef99;
aud[14202]=16'hefae;
aud[14203]=16'hefc2;
aud[14204]=16'hefd7;
aud[14205]=16'hefec;
aud[14206]=16'hf001;
aud[14207]=16'hf015;
aud[14208]=16'hf02a;
aud[14209]=16'hf03f;
aud[14210]=16'hf054;
aud[14211]=16'hf069;
aud[14212]=16'hf07d;
aud[14213]=16'hf092;
aud[14214]=16'hf0a7;
aud[14215]=16'hf0bc;
aud[14216]=16'hf0d1;
aud[14217]=16'hf0e6;
aud[14218]=16'hf0fa;
aud[14219]=16'hf10f;
aud[14220]=16'hf124;
aud[14221]=16'hf139;
aud[14222]=16'hf14e;
aud[14223]=16'hf163;
aud[14224]=16'hf178;
aud[14225]=16'hf18c;
aud[14226]=16'hf1a1;
aud[14227]=16'hf1b6;
aud[14228]=16'hf1cb;
aud[14229]=16'hf1e0;
aud[14230]=16'hf1f5;
aud[14231]=16'hf20a;
aud[14232]=16'hf21f;
aud[14233]=16'hf234;
aud[14234]=16'hf249;
aud[14235]=16'hf25e;
aud[14236]=16'hf273;
aud[14237]=16'hf288;
aud[14238]=16'hf29d;
aud[14239]=16'hf2b2;
aud[14240]=16'hf2c7;
aud[14241]=16'hf2dc;
aud[14242]=16'hf2f1;
aud[14243]=16'hf306;
aud[14244]=16'hf31b;
aud[14245]=16'hf330;
aud[14246]=16'hf345;
aud[14247]=16'hf35a;
aud[14248]=16'hf36f;
aud[14249]=16'hf384;
aud[14250]=16'hf399;
aud[14251]=16'hf3ae;
aud[14252]=16'hf3c3;
aud[14253]=16'hf3d8;
aud[14254]=16'hf3ed;
aud[14255]=16'hf402;
aud[14256]=16'hf417;
aud[14257]=16'hf42c;
aud[14258]=16'hf441;
aud[14259]=16'hf456;
aud[14260]=16'hf46b;
aud[14261]=16'hf480;
aud[14262]=16'hf496;
aud[14263]=16'hf4ab;
aud[14264]=16'hf4c0;
aud[14265]=16'hf4d5;
aud[14266]=16'hf4ea;
aud[14267]=16'hf4ff;
aud[14268]=16'hf514;
aud[14269]=16'hf529;
aud[14270]=16'hf53f;
aud[14271]=16'hf554;
aud[14272]=16'hf569;
aud[14273]=16'hf57e;
aud[14274]=16'hf593;
aud[14275]=16'hf5a8;
aud[14276]=16'hf5bd;
aud[14277]=16'hf5d3;
aud[14278]=16'hf5e8;
aud[14279]=16'hf5fd;
aud[14280]=16'hf612;
aud[14281]=16'hf627;
aud[14282]=16'hf63d;
aud[14283]=16'hf652;
aud[14284]=16'hf667;
aud[14285]=16'hf67c;
aud[14286]=16'hf691;
aud[14287]=16'hf6a7;
aud[14288]=16'hf6bc;
aud[14289]=16'hf6d1;
aud[14290]=16'hf6e6;
aud[14291]=16'hf6fb;
aud[14292]=16'hf711;
aud[14293]=16'hf726;
aud[14294]=16'hf73b;
aud[14295]=16'hf750;
aud[14296]=16'hf766;
aud[14297]=16'hf77b;
aud[14298]=16'hf790;
aud[14299]=16'hf7a5;
aud[14300]=16'hf7bb;
aud[14301]=16'hf7d0;
aud[14302]=16'hf7e5;
aud[14303]=16'hf7fb;
aud[14304]=16'hf810;
aud[14305]=16'hf825;
aud[14306]=16'hf83a;
aud[14307]=16'hf850;
aud[14308]=16'hf865;
aud[14309]=16'hf87a;
aud[14310]=16'hf890;
aud[14311]=16'hf8a5;
aud[14312]=16'hf8ba;
aud[14313]=16'hf8cf;
aud[14314]=16'hf8e5;
aud[14315]=16'hf8fa;
aud[14316]=16'hf90f;
aud[14317]=16'hf925;
aud[14318]=16'hf93a;
aud[14319]=16'hf94f;
aud[14320]=16'hf965;
aud[14321]=16'hf97a;
aud[14322]=16'hf98f;
aud[14323]=16'hf9a5;
aud[14324]=16'hf9ba;
aud[14325]=16'hf9cf;
aud[14326]=16'hf9e5;
aud[14327]=16'hf9fa;
aud[14328]=16'hfa0f;
aud[14329]=16'hfa25;
aud[14330]=16'hfa3a;
aud[14331]=16'hfa50;
aud[14332]=16'hfa65;
aud[14333]=16'hfa7a;
aud[14334]=16'hfa90;
aud[14335]=16'hfaa5;
aud[14336]=16'hfaba;
aud[14337]=16'hfad0;
aud[14338]=16'hfae5;
aud[14339]=16'hfafb;
aud[14340]=16'hfb10;
aud[14341]=16'hfb25;
aud[14342]=16'hfb3b;
aud[14343]=16'hfb50;
aud[14344]=16'hfb65;
aud[14345]=16'hfb7b;
aud[14346]=16'hfb90;
aud[14347]=16'hfba6;
aud[14348]=16'hfbbb;
aud[14349]=16'hfbd0;
aud[14350]=16'hfbe6;
aud[14351]=16'hfbfb;
aud[14352]=16'hfc11;
aud[14353]=16'hfc26;
aud[14354]=16'hfc3b;
aud[14355]=16'hfc51;
aud[14356]=16'hfc66;
aud[14357]=16'hfc7c;
aud[14358]=16'hfc91;
aud[14359]=16'hfca7;
aud[14360]=16'hfcbc;
aud[14361]=16'hfcd1;
aud[14362]=16'hfce7;
aud[14363]=16'hfcfc;
aud[14364]=16'hfd12;
aud[14365]=16'hfd27;
aud[14366]=16'hfd3c;
aud[14367]=16'hfd52;
aud[14368]=16'hfd67;
aud[14369]=16'hfd7d;
aud[14370]=16'hfd92;
aud[14371]=16'hfda8;
aud[14372]=16'hfdbd;
aud[14373]=16'hfdd2;
aud[14374]=16'hfde8;
aud[14375]=16'hfdfd;
aud[14376]=16'hfe13;
aud[14377]=16'hfe28;
aud[14378]=16'hfe3e;
aud[14379]=16'hfe53;
aud[14380]=16'hfe69;
aud[14381]=16'hfe7e;
aud[14382]=16'hfe93;
aud[14383]=16'hfea9;
aud[14384]=16'hfebe;
aud[14385]=16'hfed4;
aud[14386]=16'hfee9;
aud[14387]=16'hfeff;
aud[14388]=16'hff14;
aud[14389]=16'hff2a;
aud[14390]=16'hff3f;
aud[14391]=16'hff54;
aud[14392]=16'hff6a;
aud[14393]=16'hff7f;
aud[14394]=16'hff95;
aud[14395]=16'hffaa;
aud[14396]=16'hffc0;
aud[14397]=16'hffd5;
aud[14398]=16'hffeb;
aud[14399]=16'h0;
aud[14400]=16'h15;
aud[14401]=16'h2b;
aud[14402]=16'h40;
aud[14403]=16'h56;
aud[14404]=16'h6b;
aud[14405]=16'h81;
aud[14406]=16'h96;
aud[14407]=16'hac;
aud[14408]=16'hc1;
aud[14409]=16'hd6;
aud[14410]=16'hec;
aud[14411]=16'h101;
aud[14412]=16'h117;
aud[14413]=16'h12c;
aud[14414]=16'h142;
aud[14415]=16'h157;
aud[14416]=16'h16d;
aud[14417]=16'h182;
aud[14418]=16'h197;
aud[14419]=16'h1ad;
aud[14420]=16'h1c2;
aud[14421]=16'h1d8;
aud[14422]=16'h1ed;
aud[14423]=16'h203;
aud[14424]=16'h218;
aud[14425]=16'h22e;
aud[14426]=16'h243;
aud[14427]=16'h258;
aud[14428]=16'h26e;
aud[14429]=16'h283;
aud[14430]=16'h299;
aud[14431]=16'h2ae;
aud[14432]=16'h2c4;
aud[14433]=16'h2d9;
aud[14434]=16'h2ee;
aud[14435]=16'h304;
aud[14436]=16'h319;
aud[14437]=16'h32f;
aud[14438]=16'h344;
aud[14439]=16'h359;
aud[14440]=16'h36f;
aud[14441]=16'h384;
aud[14442]=16'h39a;
aud[14443]=16'h3af;
aud[14444]=16'h3c5;
aud[14445]=16'h3da;
aud[14446]=16'h3ef;
aud[14447]=16'h405;
aud[14448]=16'h41a;
aud[14449]=16'h430;
aud[14450]=16'h445;
aud[14451]=16'h45a;
aud[14452]=16'h470;
aud[14453]=16'h485;
aud[14454]=16'h49b;
aud[14455]=16'h4b0;
aud[14456]=16'h4c5;
aud[14457]=16'h4db;
aud[14458]=16'h4f0;
aud[14459]=16'h505;
aud[14460]=16'h51b;
aud[14461]=16'h530;
aud[14462]=16'h546;
aud[14463]=16'h55b;
aud[14464]=16'h570;
aud[14465]=16'h586;
aud[14466]=16'h59b;
aud[14467]=16'h5b0;
aud[14468]=16'h5c6;
aud[14469]=16'h5db;
aud[14470]=16'h5f1;
aud[14471]=16'h606;
aud[14472]=16'h61b;
aud[14473]=16'h631;
aud[14474]=16'h646;
aud[14475]=16'h65b;
aud[14476]=16'h671;
aud[14477]=16'h686;
aud[14478]=16'h69b;
aud[14479]=16'h6b1;
aud[14480]=16'h6c6;
aud[14481]=16'h6db;
aud[14482]=16'h6f1;
aud[14483]=16'h706;
aud[14484]=16'h71b;
aud[14485]=16'h731;
aud[14486]=16'h746;
aud[14487]=16'h75b;
aud[14488]=16'h770;
aud[14489]=16'h786;
aud[14490]=16'h79b;
aud[14491]=16'h7b0;
aud[14492]=16'h7c6;
aud[14493]=16'h7db;
aud[14494]=16'h7f0;
aud[14495]=16'h805;
aud[14496]=16'h81b;
aud[14497]=16'h830;
aud[14498]=16'h845;
aud[14499]=16'h85b;
aud[14500]=16'h870;
aud[14501]=16'h885;
aud[14502]=16'h89a;
aud[14503]=16'h8b0;
aud[14504]=16'h8c5;
aud[14505]=16'h8da;
aud[14506]=16'h8ef;
aud[14507]=16'h905;
aud[14508]=16'h91a;
aud[14509]=16'h92f;
aud[14510]=16'h944;
aud[14511]=16'h959;
aud[14512]=16'h96f;
aud[14513]=16'h984;
aud[14514]=16'h999;
aud[14515]=16'h9ae;
aud[14516]=16'h9c3;
aud[14517]=16'h9d9;
aud[14518]=16'h9ee;
aud[14519]=16'ha03;
aud[14520]=16'ha18;
aud[14521]=16'ha2d;
aud[14522]=16'ha43;
aud[14523]=16'ha58;
aud[14524]=16'ha6d;
aud[14525]=16'ha82;
aud[14526]=16'ha97;
aud[14527]=16'haac;
aud[14528]=16'hac1;
aud[14529]=16'had7;
aud[14530]=16'haec;
aud[14531]=16'hb01;
aud[14532]=16'hb16;
aud[14533]=16'hb2b;
aud[14534]=16'hb40;
aud[14535]=16'hb55;
aud[14536]=16'hb6a;
aud[14537]=16'hb80;
aud[14538]=16'hb95;
aud[14539]=16'hbaa;
aud[14540]=16'hbbf;
aud[14541]=16'hbd4;
aud[14542]=16'hbe9;
aud[14543]=16'hbfe;
aud[14544]=16'hc13;
aud[14545]=16'hc28;
aud[14546]=16'hc3d;
aud[14547]=16'hc52;
aud[14548]=16'hc67;
aud[14549]=16'hc7c;
aud[14550]=16'hc91;
aud[14551]=16'hca6;
aud[14552]=16'hcbb;
aud[14553]=16'hcd0;
aud[14554]=16'hce5;
aud[14555]=16'hcfa;
aud[14556]=16'hd0f;
aud[14557]=16'hd24;
aud[14558]=16'hd39;
aud[14559]=16'hd4e;
aud[14560]=16'hd63;
aud[14561]=16'hd78;
aud[14562]=16'hd8d;
aud[14563]=16'hda2;
aud[14564]=16'hdb7;
aud[14565]=16'hdcc;
aud[14566]=16'hde1;
aud[14567]=16'hdf6;
aud[14568]=16'he0b;
aud[14569]=16'he20;
aud[14570]=16'he35;
aud[14571]=16'he4a;
aud[14572]=16'he5f;
aud[14573]=16'he74;
aud[14574]=16'he88;
aud[14575]=16'he9d;
aud[14576]=16'heb2;
aud[14577]=16'hec7;
aud[14578]=16'hedc;
aud[14579]=16'hef1;
aud[14580]=16'hf06;
aud[14581]=16'hf1a;
aud[14582]=16'hf2f;
aud[14583]=16'hf44;
aud[14584]=16'hf59;
aud[14585]=16'hf6e;
aud[14586]=16'hf83;
aud[14587]=16'hf97;
aud[14588]=16'hfac;
aud[14589]=16'hfc1;
aud[14590]=16'hfd6;
aud[14591]=16'hfeb;
aud[14592]=16'hfff;
aud[14593]=16'h1014;
aud[14594]=16'h1029;
aud[14595]=16'h103e;
aud[14596]=16'h1052;
aud[14597]=16'h1067;
aud[14598]=16'h107c;
aud[14599]=16'h1090;
aud[14600]=16'h10a5;
aud[14601]=16'h10ba;
aud[14602]=16'h10cf;
aud[14603]=16'h10e3;
aud[14604]=16'h10f8;
aud[14605]=16'h110d;
aud[14606]=16'h1121;
aud[14607]=16'h1136;
aud[14608]=16'h114b;
aud[14609]=16'h115f;
aud[14610]=16'h1174;
aud[14611]=16'h1189;
aud[14612]=16'h119d;
aud[14613]=16'h11b2;
aud[14614]=16'h11c6;
aud[14615]=16'h11db;
aud[14616]=16'h11f0;
aud[14617]=16'h1204;
aud[14618]=16'h1219;
aud[14619]=16'h122d;
aud[14620]=16'h1242;
aud[14621]=16'h1256;
aud[14622]=16'h126b;
aud[14623]=16'h127f;
aud[14624]=16'h1294;
aud[14625]=16'h12a9;
aud[14626]=16'h12bd;
aud[14627]=16'h12d2;
aud[14628]=16'h12e6;
aud[14629]=16'h12fb;
aud[14630]=16'h130f;
aud[14631]=16'h1323;
aud[14632]=16'h1338;
aud[14633]=16'h134c;
aud[14634]=16'h1361;
aud[14635]=16'h1375;
aud[14636]=16'h138a;
aud[14637]=16'h139e;
aud[14638]=16'h13b3;
aud[14639]=16'h13c7;
aud[14640]=16'h13db;
aud[14641]=16'h13f0;
aud[14642]=16'h1404;
aud[14643]=16'h1418;
aud[14644]=16'h142d;
aud[14645]=16'h1441;
aud[14646]=16'h1455;
aud[14647]=16'h146a;
aud[14648]=16'h147e;
aud[14649]=16'h1492;
aud[14650]=16'h14a7;
aud[14651]=16'h14bb;
aud[14652]=16'h14cf;
aud[14653]=16'h14e4;
aud[14654]=16'h14f8;
aud[14655]=16'h150c;
aud[14656]=16'h1520;
aud[14657]=16'h1535;
aud[14658]=16'h1549;
aud[14659]=16'h155d;
aud[14660]=16'h1571;
aud[14661]=16'h1586;
aud[14662]=16'h159a;
aud[14663]=16'h15ae;
aud[14664]=16'h15c2;
aud[14665]=16'h15d6;
aud[14666]=16'h15ea;
aud[14667]=16'h15ff;
aud[14668]=16'h1613;
aud[14669]=16'h1627;
aud[14670]=16'h163b;
aud[14671]=16'h164f;
aud[14672]=16'h1663;
aud[14673]=16'h1677;
aud[14674]=16'h168b;
aud[14675]=16'h169f;
aud[14676]=16'h16b3;
aud[14677]=16'h16c7;
aud[14678]=16'h16db;
aud[14679]=16'h16f0;
aud[14680]=16'h1704;
aud[14681]=16'h1718;
aud[14682]=16'h172c;
aud[14683]=16'h1740;
aud[14684]=16'h1753;
aud[14685]=16'h1767;
aud[14686]=16'h177b;
aud[14687]=16'h178f;
aud[14688]=16'h17a3;
aud[14689]=16'h17b7;
aud[14690]=16'h17cb;
aud[14691]=16'h17df;
aud[14692]=16'h17f3;
aud[14693]=16'h1807;
aud[14694]=16'h181b;
aud[14695]=16'h182f;
aud[14696]=16'h1842;
aud[14697]=16'h1856;
aud[14698]=16'h186a;
aud[14699]=16'h187e;
aud[14700]=16'h1892;
aud[14701]=16'h18a5;
aud[14702]=16'h18b9;
aud[14703]=16'h18cd;
aud[14704]=16'h18e1;
aud[14705]=16'h18f5;
aud[14706]=16'h1908;
aud[14707]=16'h191c;
aud[14708]=16'h1930;
aud[14709]=16'h1943;
aud[14710]=16'h1957;
aud[14711]=16'h196b;
aud[14712]=16'h197f;
aud[14713]=16'h1992;
aud[14714]=16'h19a6;
aud[14715]=16'h19ba;
aud[14716]=16'h19cd;
aud[14717]=16'h19e1;
aud[14718]=16'h19f4;
aud[14719]=16'h1a08;
aud[14720]=16'h1a1c;
aud[14721]=16'h1a2f;
aud[14722]=16'h1a43;
aud[14723]=16'h1a56;
aud[14724]=16'h1a6a;
aud[14725]=16'h1a7d;
aud[14726]=16'h1a91;
aud[14727]=16'h1aa4;
aud[14728]=16'h1ab8;
aud[14729]=16'h1acb;
aud[14730]=16'h1adf;
aud[14731]=16'h1af2;
aud[14732]=16'h1b06;
aud[14733]=16'h1b19;
aud[14734]=16'h1b2d;
aud[14735]=16'h1b40;
aud[14736]=16'h1b53;
aud[14737]=16'h1b67;
aud[14738]=16'h1b7a;
aud[14739]=16'h1b8d;
aud[14740]=16'h1ba1;
aud[14741]=16'h1bb4;
aud[14742]=16'h1bc8;
aud[14743]=16'h1bdb;
aud[14744]=16'h1bee;
aud[14745]=16'h1c01;
aud[14746]=16'h1c15;
aud[14747]=16'h1c28;
aud[14748]=16'h1c3b;
aud[14749]=16'h1c4e;
aud[14750]=16'h1c62;
aud[14751]=16'h1c75;
aud[14752]=16'h1c88;
aud[14753]=16'h1c9b;
aud[14754]=16'h1cae;
aud[14755]=16'h1cc2;
aud[14756]=16'h1cd5;
aud[14757]=16'h1ce8;
aud[14758]=16'h1cfb;
aud[14759]=16'h1d0e;
aud[14760]=16'h1d21;
aud[14761]=16'h1d34;
aud[14762]=16'h1d47;
aud[14763]=16'h1d5b;
aud[14764]=16'h1d6e;
aud[14765]=16'h1d81;
aud[14766]=16'h1d94;
aud[14767]=16'h1da7;
aud[14768]=16'h1dba;
aud[14769]=16'h1dcd;
aud[14770]=16'h1de0;
aud[14771]=16'h1df3;
aud[14772]=16'h1e06;
aud[14773]=16'h1e18;
aud[14774]=16'h1e2b;
aud[14775]=16'h1e3e;
aud[14776]=16'h1e51;
aud[14777]=16'h1e64;
aud[14778]=16'h1e77;
aud[14779]=16'h1e8a;
aud[14780]=16'h1e9d;
aud[14781]=16'h1eaf;
aud[14782]=16'h1ec2;
aud[14783]=16'h1ed5;
aud[14784]=16'h1ee8;
aud[14785]=16'h1efb;
aud[14786]=16'h1f0d;
aud[14787]=16'h1f20;
aud[14788]=16'h1f33;
aud[14789]=16'h1f46;
aud[14790]=16'h1f58;
aud[14791]=16'h1f6b;
aud[14792]=16'h1f7e;
aud[14793]=16'h1f90;
aud[14794]=16'h1fa3;
aud[14795]=16'h1fb6;
aud[14796]=16'h1fc8;
aud[14797]=16'h1fdb;
aud[14798]=16'h1fed;
aud[14799]=16'h2000;
aud[14800]=16'h2013;
aud[14801]=16'h2025;
aud[14802]=16'h2038;
aud[14803]=16'h204a;
aud[14804]=16'h205d;
aud[14805]=16'h206f;
aud[14806]=16'h2082;
aud[14807]=16'h2094;
aud[14808]=16'h20a7;
aud[14809]=16'h20b9;
aud[14810]=16'h20cb;
aud[14811]=16'h20de;
aud[14812]=16'h20f0;
aud[14813]=16'h2103;
aud[14814]=16'h2115;
aud[14815]=16'h2127;
aud[14816]=16'h213a;
aud[14817]=16'h214c;
aud[14818]=16'h215e;
aud[14819]=16'h2171;
aud[14820]=16'h2183;
aud[14821]=16'h2195;
aud[14822]=16'h21a7;
aud[14823]=16'h21ba;
aud[14824]=16'h21cc;
aud[14825]=16'h21de;
aud[14826]=16'h21f0;
aud[14827]=16'h2202;
aud[14828]=16'h2215;
aud[14829]=16'h2227;
aud[14830]=16'h2239;
aud[14831]=16'h224b;
aud[14832]=16'h225d;
aud[14833]=16'h226f;
aud[14834]=16'h2281;
aud[14835]=16'h2293;
aud[14836]=16'h22a5;
aud[14837]=16'h22b7;
aud[14838]=16'h22c9;
aud[14839]=16'h22db;
aud[14840]=16'h22ed;
aud[14841]=16'h22ff;
aud[14842]=16'h2311;
aud[14843]=16'h2323;
aud[14844]=16'h2335;
aud[14845]=16'h2347;
aud[14846]=16'h2359;
aud[14847]=16'h236b;
aud[14848]=16'h237d;
aud[14849]=16'h238e;
aud[14850]=16'h23a0;
aud[14851]=16'h23b2;
aud[14852]=16'h23c4;
aud[14853]=16'h23d6;
aud[14854]=16'h23e7;
aud[14855]=16'h23f9;
aud[14856]=16'h240b;
aud[14857]=16'h241d;
aud[14858]=16'h242e;
aud[14859]=16'h2440;
aud[14860]=16'h2452;
aud[14861]=16'h2463;
aud[14862]=16'h2475;
aud[14863]=16'h2487;
aud[14864]=16'h2498;
aud[14865]=16'h24aa;
aud[14866]=16'h24bb;
aud[14867]=16'h24cd;
aud[14868]=16'h24de;
aud[14869]=16'h24f0;
aud[14870]=16'h2501;
aud[14871]=16'h2513;
aud[14872]=16'h2524;
aud[14873]=16'h2536;
aud[14874]=16'h2547;
aud[14875]=16'h2559;
aud[14876]=16'h256a;
aud[14877]=16'h257c;
aud[14878]=16'h258d;
aud[14879]=16'h259e;
aud[14880]=16'h25b0;
aud[14881]=16'h25c1;
aud[14882]=16'h25d2;
aud[14883]=16'h25e4;
aud[14884]=16'h25f5;
aud[14885]=16'h2606;
aud[14886]=16'h2617;
aud[14887]=16'h2629;
aud[14888]=16'h263a;
aud[14889]=16'h264b;
aud[14890]=16'h265c;
aud[14891]=16'h266d;
aud[14892]=16'h267e;
aud[14893]=16'h2690;
aud[14894]=16'h26a1;
aud[14895]=16'h26b2;
aud[14896]=16'h26c3;
aud[14897]=16'h26d4;
aud[14898]=16'h26e5;
aud[14899]=16'h26f6;
aud[14900]=16'h2707;
aud[14901]=16'h2718;
aud[14902]=16'h2729;
aud[14903]=16'h273a;
aud[14904]=16'h274b;
aud[14905]=16'h275c;
aud[14906]=16'h276d;
aud[14907]=16'h277e;
aud[14908]=16'h278e;
aud[14909]=16'h279f;
aud[14910]=16'h27b0;
aud[14911]=16'h27c1;
aud[14912]=16'h27d2;
aud[14913]=16'h27e2;
aud[14914]=16'h27f3;
aud[14915]=16'h2804;
aud[14916]=16'h2815;
aud[14917]=16'h2825;
aud[14918]=16'h2836;
aud[14919]=16'h2847;
aud[14920]=16'h2857;
aud[14921]=16'h2868;
aud[14922]=16'h2879;
aud[14923]=16'h2889;
aud[14924]=16'h289a;
aud[14925]=16'h28aa;
aud[14926]=16'h28bb;
aud[14927]=16'h28cc;
aud[14928]=16'h28dc;
aud[14929]=16'h28ed;
aud[14930]=16'h28fd;
aud[14931]=16'h290e;
aud[14932]=16'h291e;
aud[14933]=16'h292e;
aud[14934]=16'h293f;
aud[14935]=16'h294f;
aud[14936]=16'h2960;
aud[14937]=16'h2970;
aud[14938]=16'h2980;
aud[14939]=16'h2991;
aud[14940]=16'h29a1;
aud[14941]=16'h29b1;
aud[14942]=16'h29c1;
aud[14943]=16'h29d2;
aud[14944]=16'h29e2;
aud[14945]=16'h29f2;
aud[14946]=16'h2a02;
aud[14947]=16'h2a12;
aud[14948]=16'h2a23;
aud[14949]=16'h2a33;
aud[14950]=16'h2a43;
aud[14951]=16'h2a53;
aud[14952]=16'h2a63;
aud[14953]=16'h2a73;
aud[14954]=16'h2a83;
aud[14955]=16'h2a93;
aud[14956]=16'h2aa3;
aud[14957]=16'h2ab3;
aud[14958]=16'h2ac3;
aud[14959]=16'h2ad3;
aud[14960]=16'h2ae3;
aud[14961]=16'h2af3;
aud[14962]=16'h2b03;
aud[14963]=16'h2b13;
aud[14964]=16'h2b22;
aud[14965]=16'h2b32;
aud[14966]=16'h2b42;
aud[14967]=16'h2b52;
aud[14968]=16'h2b62;
aud[14969]=16'h2b71;
aud[14970]=16'h2b81;
aud[14971]=16'h2b91;
aud[14972]=16'h2ba1;
aud[14973]=16'h2bb0;
aud[14974]=16'h2bc0;
aud[14975]=16'h2bd0;
aud[14976]=16'h2bdf;
aud[14977]=16'h2bef;
aud[14978]=16'h2bfe;
aud[14979]=16'h2c0e;
aud[14980]=16'h2c1e;
aud[14981]=16'h2c2d;
aud[14982]=16'h2c3d;
aud[14983]=16'h2c4c;
aud[14984]=16'h2c5c;
aud[14985]=16'h2c6b;
aud[14986]=16'h2c7a;
aud[14987]=16'h2c8a;
aud[14988]=16'h2c99;
aud[14989]=16'h2ca9;
aud[14990]=16'h2cb8;
aud[14991]=16'h2cc7;
aud[14992]=16'h2cd7;
aud[14993]=16'h2ce6;
aud[14994]=16'h2cf5;
aud[14995]=16'h2d04;
aud[14996]=16'h2d14;
aud[14997]=16'h2d23;
aud[14998]=16'h2d32;
aud[14999]=16'h2d41;
aud[15000]=16'h2d50;
aud[15001]=16'h2d60;
aud[15002]=16'h2d6f;
aud[15003]=16'h2d7e;
aud[15004]=16'h2d8d;
aud[15005]=16'h2d9c;
aud[15006]=16'h2dab;
aud[15007]=16'h2dba;
aud[15008]=16'h2dc9;
aud[15009]=16'h2dd8;
aud[15010]=16'h2de7;
aud[15011]=16'h2df6;
aud[15012]=16'h2e05;
aud[15013]=16'h2e14;
aud[15014]=16'h2e22;
aud[15015]=16'h2e31;
aud[15016]=16'h2e40;
aud[15017]=16'h2e4f;
aud[15018]=16'h2e5e;
aud[15019]=16'h2e6d;
aud[15020]=16'h2e7b;
aud[15021]=16'h2e8a;
aud[15022]=16'h2e99;
aud[15023]=16'h2ea7;
aud[15024]=16'h2eb6;
aud[15025]=16'h2ec5;
aud[15026]=16'h2ed3;
aud[15027]=16'h2ee2;
aud[15028]=16'h2ef1;
aud[15029]=16'h2eff;
aud[15030]=16'h2f0e;
aud[15031]=16'h2f1c;
aud[15032]=16'h2f2b;
aud[15033]=16'h2f39;
aud[15034]=16'h2f48;
aud[15035]=16'h2f56;
aud[15036]=16'h2f65;
aud[15037]=16'h2f73;
aud[15038]=16'h2f81;
aud[15039]=16'h2f90;
aud[15040]=16'h2f9e;
aud[15041]=16'h2fac;
aud[15042]=16'h2fbb;
aud[15043]=16'h2fc9;
aud[15044]=16'h2fd7;
aud[15045]=16'h2fe5;
aud[15046]=16'h2ff4;
aud[15047]=16'h3002;
aud[15048]=16'h3010;
aud[15049]=16'h301e;
aud[15050]=16'h302c;
aud[15051]=16'h303a;
aud[15052]=16'h3048;
aud[15053]=16'h3057;
aud[15054]=16'h3065;
aud[15055]=16'h3073;
aud[15056]=16'h3081;
aud[15057]=16'h308f;
aud[15058]=16'h309d;
aud[15059]=16'h30aa;
aud[15060]=16'h30b8;
aud[15061]=16'h30c6;
aud[15062]=16'h30d4;
aud[15063]=16'h30e2;
aud[15064]=16'h30f0;
aud[15065]=16'h30fe;
aud[15066]=16'h310b;
aud[15067]=16'h3119;
aud[15068]=16'h3127;
aud[15069]=16'h3135;
aud[15070]=16'h3142;
aud[15071]=16'h3150;
aud[15072]=16'h315e;
aud[15073]=16'h316b;
aud[15074]=16'h3179;
aud[15075]=16'h3187;
aud[15076]=16'h3194;
aud[15077]=16'h31a2;
aud[15078]=16'h31af;
aud[15079]=16'h31bd;
aud[15080]=16'h31ca;
aud[15081]=16'h31d8;
aud[15082]=16'h31e5;
aud[15083]=16'h31f3;
aud[15084]=16'h3200;
aud[15085]=16'h320d;
aud[15086]=16'h321b;
aud[15087]=16'h3228;
aud[15088]=16'h3235;
aud[15089]=16'h3243;
aud[15090]=16'h3250;
aud[15091]=16'h325d;
aud[15092]=16'h326a;
aud[15093]=16'h3278;
aud[15094]=16'h3285;
aud[15095]=16'h3292;
aud[15096]=16'h329f;
aud[15097]=16'h32ac;
aud[15098]=16'h32b9;
aud[15099]=16'h32c6;
aud[15100]=16'h32d3;
aud[15101]=16'h32e0;
aud[15102]=16'h32ed;
aud[15103]=16'h32fa;
aud[15104]=16'h3307;
aud[15105]=16'h3314;
aud[15106]=16'h3321;
aud[15107]=16'h332e;
aud[15108]=16'h333b;
aud[15109]=16'h3348;
aud[15110]=16'h3355;
aud[15111]=16'h3361;
aud[15112]=16'h336e;
aud[15113]=16'h337b;
aud[15114]=16'h3388;
aud[15115]=16'h3394;
aud[15116]=16'h33a1;
aud[15117]=16'h33ae;
aud[15118]=16'h33ba;
aud[15119]=16'h33c7;
aud[15120]=16'h33d4;
aud[15121]=16'h33e0;
aud[15122]=16'h33ed;
aud[15123]=16'h33f9;
aud[15124]=16'h3406;
aud[15125]=16'h3412;
aud[15126]=16'h341f;
aud[15127]=16'h342b;
aud[15128]=16'h3437;
aud[15129]=16'h3444;
aud[15130]=16'h3450;
aud[15131]=16'h345d;
aud[15132]=16'h3469;
aud[15133]=16'h3475;
aud[15134]=16'h3481;
aud[15135]=16'h348e;
aud[15136]=16'h349a;
aud[15137]=16'h34a6;
aud[15138]=16'h34b2;
aud[15139]=16'h34be;
aud[15140]=16'h34cb;
aud[15141]=16'h34d7;
aud[15142]=16'h34e3;
aud[15143]=16'h34ef;
aud[15144]=16'h34fb;
aud[15145]=16'h3507;
aud[15146]=16'h3513;
aud[15147]=16'h351f;
aud[15148]=16'h352b;
aud[15149]=16'h3537;
aud[15150]=16'h3543;
aud[15151]=16'h354f;
aud[15152]=16'h355a;
aud[15153]=16'h3566;
aud[15154]=16'h3572;
aud[15155]=16'h357e;
aud[15156]=16'h358a;
aud[15157]=16'h3595;
aud[15158]=16'h35a1;
aud[15159]=16'h35ad;
aud[15160]=16'h35b8;
aud[15161]=16'h35c4;
aud[15162]=16'h35d0;
aud[15163]=16'h35db;
aud[15164]=16'h35e7;
aud[15165]=16'h35f2;
aud[15166]=16'h35fe;
aud[15167]=16'h3609;
aud[15168]=16'h3615;
aud[15169]=16'h3620;
aud[15170]=16'h362c;
aud[15171]=16'h3637;
aud[15172]=16'h3643;
aud[15173]=16'h364e;
aud[15174]=16'h3659;
aud[15175]=16'h3665;
aud[15176]=16'h3670;
aud[15177]=16'h367b;
aud[15178]=16'h3686;
aud[15179]=16'h3692;
aud[15180]=16'h369d;
aud[15181]=16'h36a8;
aud[15182]=16'h36b3;
aud[15183]=16'h36be;
aud[15184]=16'h36c9;
aud[15185]=16'h36d4;
aud[15186]=16'h36e0;
aud[15187]=16'h36eb;
aud[15188]=16'h36f6;
aud[15189]=16'h3701;
aud[15190]=16'h370b;
aud[15191]=16'h3716;
aud[15192]=16'h3721;
aud[15193]=16'h372c;
aud[15194]=16'h3737;
aud[15195]=16'h3742;
aud[15196]=16'h374d;
aud[15197]=16'h3757;
aud[15198]=16'h3762;
aud[15199]=16'h376d;
aud[15200]=16'h3778;
aud[15201]=16'h3782;
aud[15202]=16'h378d;
aud[15203]=16'h3798;
aud[15204]=16'h37a2;
aud[15205]=16'h37ad;
aud[15206]=16'h37b7;
aud[15207]=16'h37c2;
aud[15208]=16'h37cc;
aud[15209]=16'h37d7;
aud[15210]=16'h37e1;
aud[15211]=16'h37ec;
aud[15212]=16'h37f6;
aud[15213]=16'h3801;
aud[15214]=16'h380b;
aud[15215]=16'h3815;
aud[15216]=16'h3820;
aud[15217]=16'h382a;
aud[15218]=16'h3834;
aud[15219]=16'h383f;
aud[15220]=16'h3849;
aud[15221]=16'h3853;
aud[15222]=16'h385d;
aud[15223]=16'h3867;
aud[15224]=16'h3871;
aud[15225]=16'h387b;
aud[15226]=16'h3886;
aud[15227]=16'h3890;
aud[15228]=16'h389a;
aud[15229]=16'h38a4;
aud[15230]=16'h38ae;
aud[15231]=16'h38b8;
aud[15232]=16'h38c1;
aud[15233]=16'h38cb;
aud[15234]=16'h38d5;
aud[15235]=16'h38df;
aud[15236]=16'h38e9;
aud[15237]=16'h38f3;
aud[15238]=16'h38fd;
aud[15239]=16'h3906;
aud[15240]=16'h3910;
aud[15241]=16'h391a;
aud[15242]=16'h3923;
aud[15243]=16'h392d;
aud[15244]=16'h3937;
aud[15245]=16'h3940;
aud[15246]=16'h394a;
aud[15247]=16'h3953;
aud[15248]=16'h395d;
aud[15249]=16'h3966;
aud[15250]=16'h3970;
aud[15251]=16'h3979;
aud[15252]=16'h3983;
aud[15253]=16'h398c;
aud[15254]=16'h3995;
aud[15255]=16'h399f;
aud[15256]=16'h39a8;
aud[15257]=16'h39b1;
aud[15258]=16'h39bb;
aud[15259]=16'h39c4;
aud[15260]=16'h39cd;
aud[15261]=16'h39d6;
aud[15262]=16'h39e0;
aud[15263]=16'h39e9;
aud[15264]=16'h39f2;
aud[15265]=16'h39fb;
aud[15266]=16'h3a04;
aud[15267]=16'h3a0d;
aud[15268]=16'h3a16;
aud[15269]=16'h3a1f;
aud[15270]=16'h3a28;
aud[15271]=16'h3a31;
aud[15272]=16'h3a3a;
aud[15273]=16'h3a43;
aud[15274]=16'h3a4c;
aud[15275]=16'h3a54;
aud[15276]=16'h3a5d;
aud[15277]=16'h3a66;
aud[15278]=16'h3a6f;
aud[15279]=16'h3a78;
aud[15280]=16'h3a80;
aud[15281]=16'h3a89;
aud[15282]=16'h3a92;
aud[15283]=16'h3a9a;
aud[15284]=16'h3aa3;
aud[15285]=16'h3aab;
aud[15286]=16'h3ab4;
aud[15287]=16'h3abc;
aud[15288]=16'h3ac5;
aud[15289]=16'h3acd;
aud[15290]=16'h3ad6;
aud[15291]=16'h3ade;
aud[15292]=16'h3ae7;
aud[15293]=16'h3aef;
aud[15294]=16'h3af7;
aud[15295]=16'h3b00;
aud[15296]=16'h3b08;
aud[15297]=16'h3b10;
aud[15298]=16'h3b19;
aud[15299]=16'h3b21;
aud[15300]=16'h3b29;
aud[15301]=16'h3b31;
aud[15302]=16'h3b39;
aud[15303]=16'h3b41;
aud[15304]=16'h3b4a;
aud[15305]=16'h3b52;
aud[15306]=16'h3b5a;
aud[15307]=16'h3b62;
aud[15308]=16'h3b6a;
aud[15309]=16'h3b72;
aud[15310]=16'h3b7a;
aud[15311]=16'h3b81;
aud[15312]=16'h3b89;
aud[15313]=16'h3b91;
aud[15314]=16'h3b99;
aud[15315]=16'h3ba1;
aud[15316]=16'h3ba9;
aud[15317]=16'h3bb0;
aud[15318]=16'h3bb8;
aud[15319]=16'h3bc0;
aud[15320]=16'h3bc7;
aud[15321]=16'h3bcf;
aud[15322]=16'h3bd7;
aud[15323]=16'h3bde;
aud[15324]=16'h3be6;
aud[15325]=16'h3bed;
aud[15326]=16'h3bf5;
aud[15327]=16'h3bfc;
aud[15328]=16'h3c04;
aud[15329]=16'h3c0b;
aud[15330]=16'h3c13;
aud[15331]=16'h3c1a;
aud[15332]=16'h3c21;
aud[15333]=16'h3c29;
aud[15334]=16'h3c30;
aud[15335]=16'h3c37;
aud[15336]=16'h3c3f;
aud[15337]=16'h3c46;
aud[15338]=16'h3c4d;
aud[15339]=16'h3c54;
aud[15340]=16'h3c5b;
aud[15341]=16'h3c63;
aud[15342]=16'h3c6a;
aud[15343]=16'h3c71;
aud[15344]=16'h3c78;
aud[15345]=16'h3c7f;
aud[15346]=16'h3c86;
aud[15347]=16'h3c8d;
aud[15348]=16'h3c94;
aud[15349]=16'h3c9b;
aud[15350]=16'h3ca1;
aud[15351]=16'h3ca8;
aud[15352]=16'h3caf;
aud[15353]=16'h3cb6;
aud[15354]=16'h3cbd;
aud[15355]=16'h3cc3;
aud[15356]=16'h3cca;
aud[15357]=16'h3cd1;
aud[15358]=16'h3cd7;
aud[15359]=16'h3cde;
aud[15360]=16'h3ce5;
aud[15361]=16'h3ceb;
aud[15362]=16'h3cf2;
aud[15363]=16'h3cf8;
aud[15364]=16'h3cff;
aud[15365]=16'h3d05;
aud[15366]=16'h3d0c;
aud[15367]=16'h3d12;
aud[15368]=16'h3d19;
aud[15369]=16'h3d1f;
aud[15370]=16'h3d25;
aud[15371]=16'h3d2c;
aud[15372]=16'h3d32;
aud[15373]=16'h3d38;
aud[15374]=16'h3d3f;
aud[15375]=16'h3d45;
aud[15376]=16'h3d4b;
aud[15377]=16'h3d51;
aud[15378]=16'h3d57;
aud[15379]=16'h3d5d;
aud[15380]=16'h3d63;
aud[15381]=16'h3d69;
aud[15382]=16'h3d6f;
aud[15383]=16'h3d75;
aud[15384]=16'h3d7b;
aud[15385]=16'h3d81;
aud[15386]=16'h3d87;
aud[15387]=16'h3d8d;
aud[15388]=16'h3d93;
aud[15389]=16'h3d99;
aud[15390]=16'h3d9f;
aud[15391]=16'h3da4;
aud[15392]=16'h3daa;
aud[15393]=16'h3db0;
aud[15394]=16'h3db6;
aud[15395]=16'h3dbb;
aud[15396]=16'h3dc1;
aud[15397]=16'h3dc7;
aud[15398]=16'h3dcc;
aud[15399]=16'h3dd2;
aud[15400]=16'h3dd7;
aud[15401]=16'h3ddd;
aud[15402]=16'h3de2;
aud[15403]=16'h3de8;
aud[15404]=16'h3ded;
aud[15405]=16'h3df3;
aud[15406]=16'h3df8;
aud[15407]=16'h3dfd;
aud[15408]=16'h3e03;
aud[15409]=16'h3e08;
aud[15410]=16'h3e0d;
aud[15411]=16'h3e12;
aud[15412]=16'h3e18;
aud[15413]=16'h3e1d;
aud[15414]=16'h3e22;
aud[15415]=16'h3e27;
aud[15416]=16'h3e2c;
aud[15417]=16'h3e31;
aud[15418]=16'h3e36;
aud[15419]=16'h3e3b;
aud[15420]=16'h3e40;
aud[15421]=16'h3e45;
aud[15422]=16'h3e4a;
aud[15423]=16'h3e4f;
aud[15424]=16'h3e54;
aud[15425]=16'h3e59;
aud[15426]=16'h3e5e;
aud[15427]=16'h3e62;
aud[15428]=16'h3e67;
aud[15429]=16'h3e6c;
aud[15430]=16'h3e71;
aud[15431]=16'h3e75;
aud[15432]=16'h3e7a;
aud[15433]=16'h3e7f;
aud[15434]=16'h3e83;
aud[15435]=16'h3e88;
aud[15436]=16'h3e8c;
aud[15437]=16'h3e91;
aud[15438]=16'h3e95;
aud[15439]=16'h3e9a;
aud[15440]=16'h3e9e;
aud[15441]=16'h3ea3;
aud[15442]=16'h3ea7;
aud[15443]=16'h3eac;
aud[15444]=16'h3eb0;
aud[15445]=16'h3eb4;
aud[15446]=16'h3eb9;
aud[15447]=16'h3ebd;
aud[15448]=16'h3ec1;
aud[15449]=16'h3ec5;
aud[15450]=16'h3ec9;
aud[15451]=16'h3ecd;
aud[15452]=16'h3ed2;
aud[15453]=16'h3ed6;
aud[15454]=16'h3eda;
aud[15455]=16'h3ede;
aud[15456]=16'h3ee2;
aud[15457]=16'h3ee6;
aud[15458]=16'h3eea;
aud[15459]=16'h3eee;
aud[15460]=16'h3ef2;
aud[15461]=16'h3ef5;
aud[15462]=16'h3ef9;
aud[15463]=16'h3efd;
aud[15464]=16'h3f01;
aud[15465]=16'h3f05;
aud[15466]=16'h3f08;
aud[15467]=16'h3f0c;
aud[15468]=16'h3f10;
aud[15469]=16'h3f13;
aud[15470]=16'h3f17;
aud[15471]=16'h3f1b;
aud[15472]=16'h3f1e;
aud[15473]=16'h3f22;
aud[15474]=16'h3f25;
aud[15475]=16'h3f29;
aud[15476]=16'h3f2c;
aud[15477]=16'h3f30;
aud[15478]=16'h3f33;
aud[15479]=16'h3f36;
aud[15480]=16'h3f3a;
aud[15481]=16'h3f3d;
aud[15482]=16'h3f40;
aud[15483]=16'h3f43;
aud[15484]=16'h3f47;
aud[15485]=16'h3f4a;
aud[15486]=16'h3f4d;
aud[15487]=16'h3f50;
aud[15488]=16'h3f53;
aud[15489]=16'h3f56;
aud[15490]=16'h3f5a;
aud[15491]=16'h3f5d;
aud[15492]=16'h3f60;
aud[15493]=16'h3f63;
aud[15494]=16'h3f65;
aud[15495]=16'h3f68;
aud[15496]=16'h3f6b;
aud[15497]=16'h3f6e;
aud[15498]=16'h3f71;
aud[15499]=16'h3f74;
aud[15500]=16'h3f77;
aud[15501]=16'h3f79;
aud[15502]=16'h3f7c;
aud[15503]=16'h3f7f;
aud[15504]=16'h3f81;
aud[15505]=16'h3f84;
aud[15506]=16'h3f87;
aud[15507]=16'h3f89;
aud[15508]=16'h3f8c;
aud[15509]=16'h3f8e;
aud[15510]=16'h3f91;
aud[15511]=16'h3f93;
aud[15512]=16'h3f96;
aud[15513]=16'h3f98;
aud[15514]=16'h3f9b;
aud[15515]=16'h3f9d;
aud[15516]=16'h3f9f;
aud[15517]=16'h3fa2;
aud[15518]=16'h3fa4;
aud[15519]=16'h3fa6;
aud[15520]=16'h3fa8;
aud[15521]=16'h3fab;
aud[15522]=16'h3fad;
aud[15523]=16'h3faf;
aud[15524]=16'h3fb1;
aud[15525]=16'h3fb3;
aud[15526]=16'h3fb5;
aud[15527]=16'h3fb7;
aud[15528]=16'h3fb9;
aud[15529]=16'h3fbb;
aud[15530]=16'h3fbd;
aud[15531]=16'h3fbf;
aud[15532]=16'h3fc1;
aud[15533]=16'h3fc3;
aud[15534]=16'h3fc5;
aud[15535]=16'h3fc7;
aud[15536]=16'h3fc8;
aud[15537]=16'h3fca;
aud[15538]=16'h3fcc;
aud[15539]=16'h3fcd;
aud[15540]=16'h3fcf;
aud[15541]=16'h3fd1;
aud[15542]=16'h3fd2;
aud[15543]=16'h3fd4;
aud[15544]=16'h3fd6;
aud[15545]=16'h3fd7;
aud[15546]=16'h3fd9;
aud[15547]=16'h3fda;
aud[15548]=16'h3fdc;
aud[15549]=16'h3fdd;
aud[15550]=16'h3fde;
aud[15551]=16'h3fe0;
aud[15552]=16'h3fe1;
aud[15553]=16'h3fe2;
aud[15554]=16'h3fe4;
aud[15555]=16'h3fe5;
aud[15556]=16'h3fe6;
aud[15557]=16'h3fe7;
aud[15558]=16'h3fe8;
aud[15559]=16'h3fea;
aud[15560]=16'h3feb;
aud[15561]=16'h3fec;
aud[15562]=16'h3fed;
aud[15563]=16'h3fee;
aud[15564]=16'h3fef;
aud[15565]=16'h3ff0;
aud[15566]=16'h3ff1;
aud[15567]=16'h3ff2;
aud[15568]=16'h3ff3;
aud[15569]=16'h3ff3;
aud[15570]=16'h3ff4;
aud[15571]=16'h3ff5;
aud[15572]=16'h3ff6;
aud[15573]=16'h3ff7;
aud[15574]=16'h3ff7;
aud[15575]=16'h3ff8;
aud[15576]=16'h3ff9;
aud[15577]=16'h3ff9;
aud[15578]=16'h3ffa;
aud[15579]=16'h3ffa;
aud[15580]=16'h3ffb;
aud[15581]=16'h3ffb;
aud[15582]=16'h3ffc;
aud[15583]=16'h3ffc;
aud[15584]=16'h3ffd;
aud[15585]=16'h3ffd;
aud[15586]=16'h3ffe;
aud[15587]=16'h3ffe;
aud[15588]=16'h3ffe;
aud[15589]=16'h3fff;
aud[15590]=16'h3fff;
aud[15591]=16'h3fff;
aud[15592]=16'h3fff;
aud[15593]=16'h3fff;
aud[15594]=16'h4000;
aud[15595]=16'h4000;
aud[15596]=16'h4000;
aud[15597]=16'h4000;
aud[15598]=16'h4000;
aud[15599]=16'h4000;
aud[15600]=16'h4000;
aud[15601]=16'h4000;
aud[15602]=16'h4000;
aud[15603]=16'h4000;
aud[15604]=16'h4000;
aud[15605]=16'h3fff;
aud[15606]=16'h3fff;
aud[15607]=16'h3fff;
aud[15608]=16'h3fff;
aud[15609]=16'h3fff;
aud[15610]=16'h3ffe;
aud[15611]=16'h3ffe;
aud[15612]=16'h3ffe;
aud[15613]=16'h3ffd;
aud[15614]=16'h3ffd;
aud[15615]=16'h3ffc;
aud[15616]=16'h3ffc;
aud[15617]=16'h3ffb;
aud[15618]=16'h3ffb;
aud[15619]=16'h3ffa;
aud[15620]=16'h3ffa;
aud[15621]=16'h3ff9;
aud[15622]=16'h3ff9;
aud[15623]=16'h3ff8;
aud[15624]=16'h3ff7;
aud[15625]=16'h3ff7;
aud[15626]=16'h3ff6;
aud[15627]=16'h3ff5;
aud[15628]=16'h3ff4;
aud[15629]=16'h3ff3;
aud[15630]=16'h3ff3;
aud[15631]=16'h3ff2;
aud[15632]=16'h3ff1;
aud[15633]=16'h3ff0;
aud[15634]=16'h3fef;
aud[15635]=16'h3fee;
aud[15636]=16'h3fed;
aud[15637]=16'h3fec;
aud[15638]=16'h3feb;
aud[15639]=16'h3fea;
aud[15640]=16'h3fe8;
aud[15641]=16'h3fe7;
aud[15642]=16'h3fe6;
aud[15643]=16'h3fe5;
aud[15644]=16'h3fe4;
aud[15645]=16'h3fe2;
aud[15646]=16'h3fe1;
aud[15647]=16'h3fe0;
aud[15648]=16'h3fde;
aud[15649]=16'h3fdd;
aud[15650]=16'h3fdc;
aud[15651]=16'h3fda;
aud[15652]=16'h3fd9;
aud[15653]=16'h3fd7;
aud[15654]=16'h3fd6;
aud[15655]=16'h3fd4;
aud[15656]=16'h3fd2;
aud[15657]=16'h3fd1;
aud[15658]=16'h3fcf;
aud[15659]=16'h3fcd;
aud[15660]=16'h3fcc;
aud[15661]=16'h3fca;
aud[15662]=16'h3fc8;
aud[15663]=16'h3fc7;
aud[15664]=16'h3fc5;
aud[15665]=16'h3fc3;
aud[15666]=16'h3fc1;
aud[15667]=16'h3fbf;
aud[15668]=16'h3fbd;
aud[15669]=16'h3fbb;
aud[15670]=16'h3fb9;
aud[15671]=16'h3fb7;
aud[15672]=16'h3fb5;
aud[15673]=16'h3fb3;
aud[15674]=16'h3fb1;
aud[15675]=16'h3faf;
aud[15676]=16'h3fad;
aud[15677]=16'h3fab;
aud[15678]=16'h3fa8;
aud[15679]=16'h3fa6;
aud[15680]=16'h3fa4;
aud[15681]=16'h3fa2;
aud[15682]=16'h3f9f;
aud[15683]=16'h3f9d;
aud[15684]=16'h3f9b;
aud[15685]=16'h3f98;
aud[15686]=16'h3f96;
aud[15687]=16'h3f93;
aud[15688]=16'h3f91;
aud[15689]=16'h3f8e;
aud[15690]=16'h3f8c;
aud[15691]=16'h3f89;
aud[15692]=16'h3f87;
aud[15693]=16'h3f84;
aud[15694]=16'h3f81;
aud[15695]=16'h3f7f;
aud[15696]=16'h3f7c;
aud[15697]=16'h3f79;
aud[15698]=16'h3f77;
aud[15699]=16'h3f74;
aud[15700]=16'h3f71;
aud[15701]=16'h3f6e;
aud[15702]=16'h3f6b;
aud[15703]=16'h3f68;
aud[15704]=16'h3f65;
aud[15705]=16'h3f63;
aud[15706]=16'h3f60;
aud[15707]=16'h3f5d;
aud[15708]=16'h3f5a;
aud[15709]=16'h3f56;
aud[15710]=16'h3f53;
aud[15711]=16'h3f50;
aud[15712]=16'h3f4d;
aud[15713]=16'h3f4a;
aud[15714]=16'h3f47;
aud[15715]=16'h3f43;
aud[15716]=16'h3f40;
aud[15717]=16'h3f3d;
aud[15718]=16'h3f3a;
aud[15719]=16'h3f36;
aud[15720]=16'h3f33;
aud[15721]=16'h3f30;
aud[15722]=16'h3f2c;
aud[15723]=16'h3f29;
aud[15724]=16'h3f25;
aud[15725]=16'h3f22;
aud[15726]=16'h3f1e;
aud[15727]=16'h3f1b;
aud[15728]=16'h3f17;
aud[15729]=16'h3f13;
aud[15730]=16'h3f10;
aud[15731]=16'h3f0c;
aud[15732]=16'h3f08;
aud[15733]=16'h3f05;
aud[15734]=16'h3f01;
aud[15735]=16'h3efd;
aud[15736]=16'h3ef9;
aud[15737]=16'h3ef5;
aud[15738]=16'h3ef2;
aud[15739]=16'h3eee;
aud[15740]=16'h3eea;
aud[15741]=16'h3ee6;
aud[15742]=16'h3ee2;
aud[15743]=16'h3ede;
aud[15744]=16'h3eda;
aud[15745]=16'h3ed6;
aud[15746]=16'h3ed2;
aud[15747]=16'h3ecd;
aud[15748]=16'h3ec9;
aud[15749]=16'h3ec5;
aud[15750]=16'h3ec1;
aud[15751]=16'h3ebd;
aud[15752]=16'h3eb9;
aud[15753]=16'h3eb4;
aud[15754]=16'h3eb0;
aud[15755]=16'h3eac;
aud[15756]=16'h3ea7;
aud[15757]=16'h3ea3;
aud[15758]=16'h3e9e;
aud[15759]=16'h3e9a;
aud[15760]=16'h3e95;
aud[15761]=16'h3e91;
aud[15762]=16'h3e8c;
aud[15763]=16'h3e88;
aud[15764]=16'h3e83;
aud[15765]=16'h3e7f;
aud[15766]=16'h3e7a;
aud[15767]=16'h3e75;
aud[15768]=16'h3e71;
aud[15769]=16'h3e6c;
aud[15770]=16'h3e67;
aud[15771]=16'h3e62;
aud[15772]=16'h3e5e;
aud[15773]=16'h3e59;
aud[15774]=16'h3e54;
aud[15775]=16'h3e4f;
aud[15776]=16'h3e4a;
aud[15777]=16'h3e45;
aud[15778]=16'h3e40;
aud[15779]=16'h3e3b;
aud[15780]=16'h3e36;
aud[15781]=16'h3e31;
aud[15782]=16'h3e2c;
aud[15783]=16'h3e27;
aud[15784]=16'h3e22;
aud[15785]=16'h3e1d;
aud[15786]=16'h3e18;
aud[15787]=16'h3e12;
aud[15788]=16'h3e0d;
aud[15789]=16'h3e08;
aud[15790]=16'h3e03;
aud[15791]=16'h3dfd;
aud[15792]=16'h3df8;
aud[15793]=16'h3df3;
aud[15794]=16'h3ded;
aud[15795]=16'h3de8;
aud[15796]=16'h3de2;
aud[15797]=16'h3ddd;
aud[15798]=16'h3dd7;
aud[15799]=16'h3dd2;
aud[15800]=16'h3dcc;
aud[15801]=16'h3dc7;
aud[15802]=16'h3dc1;
aud[15803]=16'h3dbb;
aud[15804]=16'h3db6;
aud[15805]=16'h3db0;
aud[15806]=16'h3daa;
aud[15807]=16'h3da4;
aud[15808]=16'h3d9f;
aud[15809]=16'h3d99;
aud[15810]=16'h3d93;
aud[15811]=16'h3d8d;
aud[15812]=16'h3d87;
aud[15813]=16'h3d81;
aud[15814]=16'h3d7b;
aud[15815]=16'h3d75;
aud[15816]=16'h3d6f;
aud[15817]=16'h3d69;
aud[15818]=16'h3d63;
aud[15819]=16'h3d5d;
aud[15820]=16'h3d57;
aud[15821]=16'h3d51;
aud[15822]=16'h3d4b;
aud[15823]=16'h3d45;
aud[15824]=16'h3d3f;
aud[15825]=16'h3d38;
aud[15826]=16'h3d32;
aud[15827]=16'h3d2c;
aud[15828]=16'h3d25;
aud[15829]=16'h3d1f;
aud[15830]=16'h3d19;
aud[15831]=16'h3d12;
aud[15832]=16'h3d0c;
aud[15833]=16'h3d05;
aud[15834]=16'h3cff;
aud[15835]=16'h3cf8;
aud[15836]=16'h3cf2;
aud[15837]=16'h3ceb;
aud[15838]=16'h3ce5;
aud[15839]=16'h3cde;
aud[15840]=16'h3cd7;
aud[15841]=16'h3cd1;
aud[15842]=16'h3cca;
aud[15843]=16'h3cc3;
aud[15844]=16'h3cbd;
aud[15845]=16'h3cb6;
aud[15846]=16'h3caf;
aud[15847]=16'h3ca8;
aud[15848]=16'h3ca1;
aud[15849]=16'h3c9b;
aud[15850]=16'h3c94;
aud[15851]=16'h3c8d;
aud[15852]=16'h3c86;
aud[15853]=16'h3c7f;
aud[15854]=16'h3c78;
aud[15855]=16'h3c71;
aud[15856]=16'h3c6a;
aud[15857]=16'h3c63;
aud[15858]=16'h3c5b;
aud[15859]=16'h3c54;
aud[15860]=16'h3c4d;
aud[15861]=16'h3c46;
aud[15862]=16'h3c3f;
aud[15863]=16'h3c37;
aud[15864]=16'h3c30;
aud[15865]=16'h3c29;
aud[15866]=16'h3c21;
aud[15867]=16'h3c1a;
aud[15868]=16'h3c13;
aud[15869]=16'h3c0b;
aud[15870]=16'h3c04;
aud[15871]=16'h3bfc;
aud[15872]=16'h3bf5;
aud[15873]=16'h3bed;
aud[15874]=16'h3be6;
aud[15875]=16'h3bde;
aud[15876]=16'h3bd7;
aud[15877]=16'h3bcf;
aud[15878]=16'h3bc7;
aud[15879]=16'h3bc0;
aud[15880]=16'h3bb8;
aud[15881]=16'h3bb0;
aud[15882]=16'h3ba9;
aud[15883]=16'h3ba1;
aud[15884]=16'h3b99;
aud[15885]=16'h3b91;
aud[15886]=16'h3b89;
aud[15887]=16'h3b81;
aud[15888]=16'h3b7a;
aud[15889]=16'h3b72;
aud[15890]=16'h3b6a;
aud[15891]=16'h3b62;
aud[15892]=16'h3b5a;
aud[15893]=16'h3b52;
aud[15894]=16'h3b4a;
aud[15895]=16'h3b41;
aud[15896]=16'h3b39;
aud[15897]=16'h3b31;
aud[15898]=16'h3b29;
aud[15899]=16'h3b21;
aud[15900]=16'h3b19;
aud[15901]=16'h3b10;
aud[15902]=16'h3b08;
aud[15903]=16'h3b00;
aud[15904]=16'h3af7;
aud[15905]=16'h3aef;
aud[15906]=16'h3ae7;
aud[15907]=16'h3ade;
aud[15908]=16'h3ad6;
aud[15909]=16'h3acd;
aud[15910]=16'h3ac5;
aud[15911]=16'h3abc;
aud[15912]=16'h3ab4;
aud[15913]=16'h3aab;
aud[15914]=16'h3aa3;
aud[15915]=16'h3a9a;
aud[15916]=16'h3a92;
aud[15917]=16'h3a89;
aud[15918]=16'h3a80;
aud[15919]=16'h3a78;
aud[15920]=16'h3a6f;
aud[15921]=16'h3a66;
aud[15922]=16'h3a5d;
aud[15923]=16'h3a54;
aud[15924]=16'h3a4c;
aud[15925]=16'h3a43;
aud[15926]=16'h3a3a;
aud[15927]=16'h3a31;
aud[15928]=16'h3a28;
aud[15929]=16'h3a1f;
aud[15930]=16'h3a16;
aud[15931]=16'h3a0d;
aud[15932]=16'h3a04;
aud[15933]=16'h39fb;
aud[15934]=16'h39f2;
aud[15935]=16'h39e9;
aud[15936]=16'h39e0;
aud[15937]=16'h39d6;
aud[15938]=16'h39cd;
aud[15939]=16'h39c4;
aud[15940]=16'h39bb;
aud[15941]=16'h39b1;
aud[15942]=16'h39a8;
aud[15943]=16'h399f;
aud[15944]=16'h3995;
aud[15945]=16'h398c;
aud[15946]=16'h3983;
aud[15947]=16'h3979;
aud[15948]=16'h3970;
aud[15949]=16'h3966;
aud[15950]=16'h395d;
aud[15951]=16'h3953;
aud[15952]=16'h394a;
aud[15953]=16'h3940;
aud[15954]=16'h3937;
aud[15955]=16'h392d;
aud[15956]=16'h3923;
aud[15957]=16'h391a;
aud[15958]=16'h3910;
aud[15959]=16'h3906;
aud[15960]=16'h38fd;
aud[15961]=16'h38f3;
aud[15962]=16'h38e9;
aud[15963]=16'h38df;
aud[15964]=16'h38d5;
aud[15965]=16'h38cb;
aud[15966]=16'h38c1;
aud[15967]=16'h38b8;
aud[15968]=16'h38ae;
aud[15969]=16'h38a4;
aud[15970]=16'h389a;
aud[15971]=16'h3890;
aud[15972]=16'h3886;
aud[15973]=16'h387b;
aud[15974]=16'h3871;
aud[15975]=16'h3867;
aud[15976]=16'h385d;
aud[15977]=16'h3853;
aud[15978]=16'h3849;
aud[15979]=16'h383f;
aud[15980]=16'h3834;
aud[15981]=16'h382a;
aud[15982]=16'h3820;
aud[15983]=16'h3815;
aud[15984]=16'h380b;
aud[15985]=16'h3801;
aud[15986]=16'h37f6;
aud[15987]=16'h37ec;
aud[15988]=16'h37e1;
aud[15989]=16'h37d7;
aud[15990]=16'h37cc;
aud[15991]=16'h37c2;
aud[15992]=16'h37b7;
aud[15993]=16'h37ad;
aud[15994]=16'h37a2;
aud[15995]=16'h3798;
aud[15996]=16'h378d;
aud[15997]=16'h3782;
aud[15998]=16'h3778;
aud[15999]=16'h376d;
aud[16000]=16'h3762;
aud[16001]=16'h3757;
aud[16002]=16'h374d;
aud[16003]=16'h3742;
aud[16004]=16'h3737;
aud[16005]=16'h372c;
aud[16006]=16'h3721;
aud[16007]=16'h3716;
aud[16008]=16'h370b;
aud[16009]=16'h3701;
aud[16010]=16'h36f6;
aud[16011]=16'h36eb;
aud[16012]=16'h36e0;
aud[16013]=16'h36d4;
aud[16014]=16'h36c9;
aud[16015]=16'h36be;
aud[16016]=16'h36b3;
aud[16017]=16'h36a8;
aud[16018]=16'h369d;
aud[16019]=16'h3692;
aud[16020]=16'h3686;
aud[16021]=16'h367b;
aud[16022]=16'h3670;
aud[16023]=16'h3665;
aud[16024]=16'h3659;
aud[16025]=16'h364e;
aud[16026]=16'h3643;
aud[16027]=16'h3637;
aud[16028]=16'h362c;
aud[16029]=16'h3620;
aud[16030]=16'h3615;
aud[16031]=16'h3609;
aud[16032]=16'h35fe;
aud[16033]=16'h35f2;
aud[16034]=16'h35e7;
aud[16035]=16'h35db;
aud[16036]=16'h35d0;
aud[16037]=16'h35c4;
aud[16038]=16'h35b8;
aud[16039]=16'h35ad;
aud[16040]=16'h35a1;
aud[16041]=16'h3595;
aud[16042]=16'h358a;
aud[16043]=16'h357e;
aud[16044]=16'h3572;
aud[16045]=16'h3566;
aud[16046]=16'h355a;
aud[16047]=16'h354f;
aud[16048]=16'h3543;
aud[16049]=16'h3537;
aud[16050]=16'h352b;
aud[16051]=16'h351f;
aud[16052]=16'h3513;
aud[16053]=16'h3507;
aud[16054]=16'h34fb;
aud[16055]=16'h34ef;
aud[16056]=16'h34e3;
aud[16057]=16'h34d7;
aud[16058]=16'h34cb;
aud[16059]=16'h34be;
aud[16060]=16'h34b2;
aud[16061]=16'h34a6;
aud[16062]=16'h349a;
aud[16063]=16'h348e;
aud[16064]=16'h3481;
aud[16065]=16'h3475;
aud[16066]=16'h3469;
aud[16067]=16'h345d;
aud[16068]=16'h3450;
aud[16069]=16'h3444;
aud[16070]=16'h3437;
aud[16071]=16'h342b;
aud[16072]=16'h341f;
aud[16073]=16'h3412;
aud[16074]=16'h3406;
aud[16075]=16'h33f9;
aud[16076]=16'h33ed;
aud[16077]=16'h33e0;
aud[16078]=16'h33d4;
aud[16079]=16'h33c7;
aud[16080]=16'h33ba;
aud[16081]=16'h33ae;
aud[16082]=16'h33a1;
aud[16083]=16'h3394;
aud[16084]=16'h3388;
aud[16085]=16'h337b;
aud[16086]=16'h336e;
aud[16087]=16'h3361;
aud[16088]=16'h3355;
aud[16089]=16'h3348;
aud[16090]=16'h333b;
aud[16091]=16'h332e;
aud[16092]=16'h3321;
aud[16093]=16'h3314;
aud[16094]=16'h3307;
aud[16095]=16'h32fa;
aud[16096]=16'h32ed;
aud[16097]=16'h32e0;
aud[16098]=16'h32d3;
aud[16099]=16'h32c6;
aud[16100]=16'h32b9;
aud[16101]=16'h32ac;
aud[16102]=16'h329f;
aud[16103]=16'h3292;
aud[16104]=16'h3285;
aud[16105]=16'h3278;
aud[16106]=16'h326a;
aud[16107]=16'h325d;
aud[16108]=16'h3250;
aud[16109]=16'h3243;
aud[16110]=16'h3235;
aud[16111]=16'h3228;
aud[16112]=16'h321b;
aud[16113]=16'h320d;
aud[16114]=16'h3200;
aud[16115]=16'h31f3;
aud[16116]=16'h31e5;
aud[16117]=16'h31d8;
aud[16118]=16'h31ca;
aud[16119]=16'h31bd;
aud[16120]=16'h31af;
aud[16121]=16'h31a2;
aud[16122]=16'h3194;
aud[16123]=16'h3187;
aud[16124]=16'h3179;
aud[16125]=16'h316b;
aud[16126]=16'h315e;
aud[16127]=16'h3150;
aud[16128]=16'h3142;
aud[16129]=16'h3135;
aud[16130]=16'h3127;
aud[16131]=16'h3119;
aud[16132]=16'h310b;
aud[16133]=16'h30fe;
aud[16134]=16'h30f0;
aud[16135]=16'h30e2;
aud[16136]=16'h30d4;
aud[16137]=16'h30c6;
aud[16138]=16'h30b8;
aud[16139]=16'h30aa;
aud[16140]=16'h309d;
aud[16141]=16'h308f;
aud[16142]=16'h3081;
aud[16143]=16'h3073;
aud[16144]=16'h3065;
aud[16145]=16'h3057;
aud[16146]=16'h3048;
aud[16147]=16'h303a;
aud[16148]=16'h302c;
aud[16149]=16'h301e;
aud[16150]=16'h3010;
aud[16151]=16'h3002;
aud[16152]=16'h2ff4;
aud[16153]=16'h2fe5;
aud[16154]=16'h2fd7;
aud[16155]=16'h2fc9;
aud[16156]=16'h2fbb;
aud[16157]=16'h2fac;
aud[16158]=16'h2f9e;
aud[16159]=16'h2f90;
aud[16160]=16'h2f81;
aud[16161]=16'h2f73;
aud[16162]=16'h2f65;
aud[16163]=16'h2f56;
aud[16164]=16'h2f48;
aud[16165]=16'h2f39;
aud[16166]=16'h2f2b;
aud[16167]=16'h2f1c;
aud[16168]=16'h2f0e;
aud[16169]=16'h2eff;
aud[16170]=16'h2ef1;
aud[16171]=16'h2ee2;
aud[16172]=16'h2ed3;
aud[16173]=16'h2ec5;
aud[16174]=16'h2eb6;
aud[16175]=16'h2ea7;
aud[16176]=16'h2e99;
aud[16177]=16'h2e8a;
aud[16178]=16'h2e7b;
aud[16179]=16'h2e6d;
aud[16180]=16'h2e5e;
aud[16181]=16'h2e4f;
aud[16182]=16'h2e40;
aud[16183]=16'h2e31;
aud[16184]=16'h2e22;
aud[16185]=16'h2e14;
aud[16186]=16'h2e05;
aud[16187]=16'h2df6;
aud[16188]=16'h2de7;
aud[16189]=16'h2dd8;
aud[16190]=16'h2dc9;
aud[16191]=16'h2dba;
aud[16192]=16'h2dab;
aud[16193]=16'h2d9c;
aud[16194]=16'h2d8d;
aud[16195]=16'h2d7e;
aud[16196]=16'h2d6f;
aud[16197]=16'h2d60;
aud[16198]=16'h2d50;
aud[16199]=16'h2d41;
aud[16200]=16'h2d32;
aud[16201]=16'h2d23;
aud[16202]=16'h2d14;
aud[16203]=16'h2d04;
aud[16204]=16'h2cf5;
aud[16205]=16'h2ce6;
aud[16206]=16'h2cd7;
aud[16207]=16'h2cc7;
aud[16208]=16'h2cb8;
aud[16209]=16'h2ca9;
aud[16210]=16'h2c99;
aud[16211]=16'h2c8a;
aud[16212]=16'h2c7a;
aud[16213]=16'h2c6b;
aud[16214]=16'h2c5c;
aud[16215]=16'h2c4c;
aud[16216]=16'h2c3d;
aud[16217]=16'h2c2d;
aud[16218]=16'h2c1e;
aud[16219]=16'h2c0e;
aud[16220]=16'h2bfe;
aud[16221]=16'h2bef;
aud[16222]=16'h2bdf;
aud[16223]=16'h2bd0;
aud[16224]=16'h2bc0;
aud[16225]=16'h2bb0;
aud[16226]=16'h2ba1;
aud[16227]=16'h2b91;
aud[16228]=16'h2b81;
aud[16229]=16'h2b71;
aud[16230]=16'h2b62;
aud[16231]=16'h2b52;
aud[16232]=16'h2b42;
aud[16233]=16'h2b32;
aud[16234]=16'h2b22;
aud[16235]=16'h2b13;
aud[16236]=16'h2b03;
aud[16237]=16'h2af3;
aud[16238]=16'h2ae3;
aud[16239]=16'h2ad3;
aud[16240]=16'h2ac3;
aud[16241]=16'h2ab3;
aud[16242]=16'h2aa3;
aud[16243]=16'h2a93;
aud[16244]=16'h2a83;
aud[16245]=16'h2a73;
aud[16246]=16'h2a63;
aud[16247]=16'h2a53;
aud[16248]=16'h2a43;
aud[16249]=16'h2a33;
aud[16250]=16'h2a23;
aud[16251]=16'h2a12;
aud[16252]=16'h2a02;
aud[16253]=16'h29f2;
aud[16254]=16'h29e2;
aud[16255]=16'h29d2;
aud[16256]=16'h29c1;
aud[16257]=16'h29b1;
aud[16258]=16'h29a1;
aud[16259]=16'h2991;
aud[16260]=16'h2980;
aud[16261]=16'h2970;
aud[16262]=16'h2960;
aud[16263]=16'h294f;
aud[16264]=16'h293f;
aud[16265]=16'h292e;
aud[16266]=16'h291e;
aud[16267]=16'h290e;
aud[16268]=16'h28fd;
aud[16269]=16'h28ed;
aud[16270]=16'h28dc;
aud[16271]=16'h28cc;
aud[16272]=16'h28bb;
aud[16273]=16'h28aa;
aud[16274]=16'h289a;
aud[16275]=16'h2889;
aud[16276]=16'h2879;
aud[16277]=16'h2868;
aud[16278]=16'h2857;
aud[16279]=16'h2847;
aud[16280]=16'h2836;
aud[16281]=16'h2825;
aud[16282]=16'h2815;
aud[16283]=16'h2804;
aud[16284]=16'h27f3;
aud[16285]=16'h27e2;
aud[16286]=16'h27d2;
aud[16287]=16'h27c1;
aud[16288]=16'h27b0;
aud[16289]=16'h279f;
aud[16290]=16'h278e;
aud[16291]=16'h277e;
aud[16292]=16'h276d;
aud[16293]=16'h275c;
aud[16294]=16'h274b;
aud[16295]=16'h273a;
aud[16296]=16'h2729;
aud[16297]=16'h2718;
aud[16298]=16'h2707;
aud[16299]=16'h26f6;
aud[16300]=16'h26e5;
aud[16301]=16'h26d4;
aud[16302]=16'h26c3;
aud[16303]=16'h26b2;
aud[16304]=16'h26a1;
aud[16305]=16'h2690;
aud[16306]=16'h267e;
aud[16307]=16'h266d;
aud[16308]=16'h265c;
aud[16309]=16'h264b;
aud[16310]=16'h263a;
aud[16311]=16'h2629;
aud[16312]=16'h2617;
aud[16313]=16'h2606;
aud[16314]=16'h25f5;
aud[16315]=16'h25e4;
aud[16316]=16'h25d2;
aud[16317]=16'h25c1;
aud[16318]=16'h25b0;
aud[16319]=16'h259e;
aud[16320]=16'h258d;
aud[16321]=16'h257c;
aud[16322]=16'h256a;
aud[16323]=16'h2559;
aud[16324]=16'h2547;
aud[16325]=16'h2536;
aud[16326]=16'h2524;
aud[16327]=16'h2513;
aud[16328]=16'h2501;
aud[16329]=16'h24f0;
aud[16330]=16'h24de;
aud[16331]=16'h24cd;
aud[16332]=16'h24bb;
aud[16333]=16'h24aa;
aud[16334]=16'h2498;
aud[16335]=16'h2487;
aud[16336]=16'h2475;
aud[16337]=16'h2463;
aud[16338]=16'h2452;
aud[16339]=16'h2440;
aud[16340]=16'h242e;
aud[16341]=16'h241d;
aud[16342]=16'h240b;
aud[16343]=16'h23f9;
aud[16344]=16'h23e7;
aud[16345]=16'h23d6;
aud[16346]=16'h23c4;
aud[16347]=16'h23b2;
aud[16348]=16'h23a0;
aud[16349]=16'h238e;
aud[16350]=16'h237d;
aud[16351]=16'h236b;
aud[16352]=16'h2359;
aud[16353]=16'h2347;
aud[16354]=16'h2335;
aud[16355]=16'h2323;
aud[16356]=16'h2311;
aud[16357]=16'h22ff;
aud[16358]=16'h22ed;
aud[16359]=16'h22db;
aud[16360]=16'h22c9;
aud[16361]=16'h22b7;
aud[16362]=16'h22a5;
aud[16363]=16'h2293;
aud[16364]=16'h2281;
aud[16365]=16'h226f;
aud[16366]=16'h225d;
aud[16367]=16'h224b;
aud[16368]=16'h2239;
aud[16369]=16'h2227;
aud[16370]=16'h2215;
aud[16371]=16'h2202;
aud[16372]=16'h21f0;
aud[16373]=16'h21de;
aud[16374]=16'h21cc;
aud[16375]=16'h21ba;
aud[16376]=16'h21a7;
aud[16377]=16'h2195;
aud[16378]=16'h2183;
aud[16379]=16'h2171;
aud[16380]=16'h215e;
aud[16381]=16'h214c;
aud[16382]=16'h213a;
aud[16383]=16'h2127;
aud[16384]=16'h2115;
aud[16385]=16'h2103;
aud[16386]=16'h20f0;
aud[16387]=16'h20de;
aud[16388]=16'h20cb;
aud[16389]=16'h20b9;
aud[16390]=16'h20a7;
aud[16391]=16'h2094;
aud[16392]=16'h2082;
aud[16393]=16'h206f;
aud[16394]=16'h205d;
aud[16395]=16'h204a;
aud[16396]=16'h2038;
aud[16397]=16'h2025;
aud[16398]=16'h2013;
aud[16399]=16'h2000;
aud[16400]=16'h1fed;
aud[16401]=16'h1fdb;
aud[16402]=16'h1fc8;
aud[16403]=16'h1fb6;
aud[16404]=16'h1fa3;
aud[16405]=16'h1f90;
aud[16406]=16'h1f7e;
aud[16407]=16'h1f6b;
aud[16408]=16'h1f58;
aud[16409]=16'h1f46;
aud[16410]=16'h1f33;
aud[16411]=16'h1f20;
aud[16412]=16'h1f0d;
aud[16413]=16'h1efb;
aud[16414]=16'h1ee8;
aud[16415]=16'h1ed5;
aud[16416]=16'h1ec2;
aud[16417]=16'h1eaf;
aud[16418]=16'h1e9d;
aud[16419]=16'h1e8a;
aud[16420]=16'h1e77;
aud[16421]=16'h1e64;
aud[16422]=16'h1e51;
aud[16423]=16'h1e3e;
aud[16424]=16'h1e2b;
aud[16425]=16'h1e18;
aud[16426]=16'h1e06;
aud[16427]=16'h1df3;
aud[16428]=16'h1de0;
aud[16429]=16'h1dcd;
aud[16430]=16'h1dba;
aud[16431]=16'h1da7;
aud[16432]=16'h1d94;
aud[16433]=16'h1d81;
aud[16434]=16'h1d6e;
aud[16435]=16'h1d5b;
aud[16436]=16'h1d47;
aud[16437]=16'h1d34;
aud[16438]=16'h1d21;
aud[16439]=16'h1d0e;
aud[16440]=16'h1cfb;
aud[16441]=16'h1ce8;
aud[16442]=16'h1cd5;
aud[16443]=16'h1cc2;
aud[16444]=16'h1cae;
aud[16445]=16'h1c9b;
aud[16446]=16'h1c88;
aud[16447]=16'h1c75;
aud[16448]=16'h1c62;
aud[16449]=16'h1c4e;
aud[16450]=16'h1c3b;
aud[16451]=16'h1c28;
aud[16452]=16'h1c15;
aud[16453]=16'h1c01;
aud[16454]=16'h1bee;
aud[16455]=16'h1bdb;
aud[16456]=16'h1bc8;
aud[16457]=16'h1bb4;
aud[16458]=16'h1ba1;
aud[16459]=16'h1b8d;
aud[16460]=16'h1b7a;
aud[16461]=16'h1b67;
aud[16462]=16'h1b53;
aud[16463]=16'h1b40;
aud[16464]=16'h1b2d;
aud[16465]=16'h1b19;
aud[16466]=16'h1b06;
aud[16467]=16'h1af2;
aud[16468]=16'h1adf;
aud[16469]=16'h1acb;
aud[16470]=16'h1ab8;
aud[16471]=16'h1aa4;
aud[16472]=16'h1a91;
aud[16473]=16'h1a7d;
aud[16474]=16'h1a6a;
aud[16475]=16'h1a56;
aud[16476]=16'h1a43;
aud[16477]=16'h1a2f;
aud[16478]=16'h1a1c;
aud[16479]=16'h1a08;
aud[16480]=16'h19f4;
aud[16481]=16'h19e1;
aud[16482]=16'h19cd;
aud[16483]=16'h19ba;
aud[16484]=16'h19a6;
aud[16485]=16'h1992;
aud[16486]=16'h197f;
aud[16487]=16'h196b;
aud[16488]=16'h1957;
aud[16489]=16'h1943;
aud[16490]=16'h1930;
aud[16491]=16'h191c;
aud[16492]=16'h1908;
aud[16493]=16'h18f5;
aud[16494]=16'h18e1;
aud[16495]=16'h18cd;
aud[16496]=16'h18b9;
aud[16497]=16'h18a5;
aud[16498]=16'h1892;
aud[16499]=16'h187e;
aud[16500]=16'h186a;
aud[16501]=16'h1856;
aud[16502]=16'h1842;
aud[16503]=16'h182f;
aud[16504]=16'h181b;
aud[16505]=16'h1807;
aud[16506]=16'h17f3;
aud[16507]=16'h17df;
aud[16508]=16'h17cb;
aud[16509]=16'h17b7;
aud[16510]=16'h17a3;
aud[16511]=16'h178f;
aud[16512]=16'h177b;
aud[16513]=16'h1767;
aud[16514]=16'h1753;
aud[16515]=16'h1740;
aud[16516]=16'h172c;
aud[16517]=16'h1718;
aud[16518]=16'h1704;
aud[16519]=16'h16f0;
aud[16520]=16'h16db;
aud[16521]=16'h16c7;
aud[16522]=16'h16b3;
aud[16523]=16'h169f;
aud[16524]=16'h168b;
aud[16525]=16'h1677;
aud[16526]=16'h1663;
aud[16527]=16'h164f;
aud[16528]=16'h163b;
aud[16529]=16'h1627;
aud[16530]=16'h1613;
aud[16531]=16'h15ff;
aud[16532]=16'h15ea;
aud[16533]=16'h15d6;
aud[16534]=16'h15c2;
aud[16535]=16'h15ae;
aud[16536]=16'h159a;
aud[16537]=16'h1586;
aud[16538]=16'h1571;
aud[16539]=16'h155d;
aud[16540]=16'h1549;
aud[16541]=16'h1535;
aud[16542]=16'h1520;
aud[16543]=16'h150c;
aud[16544]=16'h14f8;
aud[16545]=16'h14e4;
aud[16546]=16'h14cf;
aud[16547]=16'h14bb;
aud[16548]=16'h14a7;
aud[16549]=16'h1492;
aud[16550]=16'h147e;
aud[16551]=16'h146a;
aud[16552]=16'h1455;
aud[16553]=16'h1441;
aud[16554]=16'h142d;
aud[16555]=16'h1418;
aud[16556]=16'h1404;
aud[16557]=16'h13f0;
aud[16558]=16'h13db;
aud[16559]=16'h13c7;
aud[16560]=16'h13b3;
aud[16561]=16'h139e;
aud[16562]=16'h138a;
aud[16563]=16'h1375;
aud[16564]=16'h1361;
aud[16565]=16'h134c;
aud[16566]=16'h1338;
aud[16567]=16'h1323;
aud[16568]=16'h130f;
aud[16569]=16'h12fb;
aud[16570]=16'h12e6;
aud[16571]=16'h12d2;
aud[16572]=16'h12bd;
aud[16573]=16'h12a9;
aud[16574]=16'h1294;
aud[16575]=16'h127f;
aud[16576]=16'h126b;
aud[16577]=16'h1256;
aud[16578]=16'h1242;
aud[16579]=16'h122d;
aud[16580]=16'h1219;
aud[16581]=16'h1204;
aud[16582]=16'h11f0;
aud[16583]=16'h11db;
aud[16584]=16'h11c6;
aud[16585]=16'h11b2;
aud[16586]=16'h119d;
aud[16587]=16'h1189;
aud[16588]=16'h1174;
aud[16589]=16'h115f;
aud[16590]=16'h114b;
aud[16591]=16'h1136;
aud[16592]=16'h1121;
aud[16593]=16'h110d;
aud[16594]=16'h10f8;
aud[16595]=16'h10e3;
aud[16596]=16'h10cf;
aud[16597]=16'h10ba;
aud[16598]=16'h10a5;
aud[16599]=16'h1090;
aud[16600]=16'h107c;
aud[16601]=16'h1067;
aud[16602]=16'h1052;
aud[16603]=16'h103e;
aud[16604]=16'h1029;
aud[16605]=16'h1014;
aud[16606]=16'hfff;
aud[16607]=16'hfeb;
aud[16608]=16'hfd6;
aud[16609]=16'hfc1;
aud[16610]=16'hfac;
aud[16611]=16'hf97;
aud[16612]=16'hf83;
aud[16613]=16'hf6e;
aud[16614]=16'hf59;
aud[16615]=16'hf44;
aud[16616]=16'hf2f;
aud[16617]=16'hf1a;
aud[16618]=16'hf06;
aud[16619]=16'hef1;
aud[16620]=16'hedc;
aud[16621]=16'hec7;
aud[16622]=16'heb2;
aud[16623]=16'he9d;
aud[16624]=16'he88;
aud[16625]=16'he74;
aud[16626]=16'he5f;
aud[16627]=16'he4a;
aud[16628]=16'he35;
aud[16629]=16'he20;
aud[16630]=16'he0b;
aud[16631]=16'hdf6;
aud[16632]=16'hde1;
aud[16633]=16'hdcc;
aud[16634]=16'hdb7;
aud[16635]=16'hda2;
aud[16636]=16'hd8d;
aud[16637]=16'hd78;
aud[16638]=16'hd63;
aud[16639]=16'hd4e;
aud[16640]=16'hd39;
aud[16641]=16'hd24;
aud[16642]=16'hd0f;
aud[16643]=16'hcfa;
aud[16644]=16'hce5;
aud[16645]=16'hcd0;
aud[16646]=16'hcbb;
aud[16647]=16'hca6;
aud[16648]=16'hc91;
aud[16649]=16'hc7c;
aud[16650]=16'hc67;
aud[16651]=16'hc52;
aud[16652]=16'hc3d;
aud[16653]=16'hc28;
aud[16654]=16'hc13;
aud[16655]=16'hbfe;
aud[16656]=16'hbe9;
aud[16657]=16'hbd4;
aud[16658]=16'hbbf;
aud[16659]=16'hbaa;
aud[16660]=16'hb95;
aud[16661]=16'hb80;
aud[16662]=16'hb6a;
aud[16663]=16'hb55;
aud[16664]=16'hb40;
aud[16665]=16'hb2b;
aud[16666]=16'hb16;
aud[16667]=16'hb01;
aud[16668]=16'haec;
aud[16669]=16'had7;
aud[16670]=16'hac1;
aud[16671]=16'haac;
aud[16672]=16'ha97;
aud[16673]=16'ha82;
aud[16674]=16'ha6d;
aud[16675]=16'ha58;
aud[16676]=16'ha43;
aud[16677]=16'ha2d;
aud[16678]=16'ha18;
aud[16679]=16'ha03;
aud[16680]=16'h9ee;
aud[16681]=16'h9d9;
aud[16682]=16'h9c3;
aud[16683]=16'h9ae;
aud[16684]=16'h999;
aud[16685]=16'h984;
aud[16686]=16'h96f;
aud[16687]=16'h959;
aud[16688]=16'h944;
aud[16689]=16'h92f;
aud[16690]=16'h91a;
aud[16691]=16'h905;
aud[16692]=16'h8ef;
aud[16693]=16'h8da;
aud[16694]=16'h8c5;
aud[16695]=16'h8b0;
aud[16696]=16'h89a;
aud[16697]=16'h885;
aud[16698]=16'h870;
aud[16699]=16'h85b;
aud[16700]=16'h845;
aud[16701]=16'h830;
aud[16702]=16'h81b;
aud[16703]=16'h805;
aud[16704]=16'h7f0;
aud[16705]=16'h7db;
aud[16706]=16'h7c6;
aud[16707]=16'h7b0;
aud[16708]=16'h79b;
aud[16709]=16'h786;
aud[16710]=16'h770;
aud[16711]=16'h75b;
aud[16712]=16'h746;
aud[16713]=16'h731;
aud[16714]=16'h71b;
aud[16715]=16'h706;
aud[16716]=16'h6f1;
aud[16717]=16'h6db;
aud[16718]=16'h6c6;
aud[16719]=16'h6b1;
aud[16720]=16'h69b;
aud[16721]=16'h686;
aud[16722]=16'h671;
aud[16723]=16'h65b;
aud[16724]=16'h646;
aud[16725]=16'h631;
aud[16726]=16'h61b;
aud[16727]=16'h606;
aud[16728]=16'h5f1;
aud[16729]=16'h5db;
aud[16730]=16'h5c6;
aud[16731]=16'h5b0;
aud[16732]=16'h59b;
aud[16733]=16'h586;
aud[16734]=16'h570;
aud[16735]=16'h55b;
aud[16736]=16'h546;
aud[16737]=16'h530;
aud[16738]=16'h51b;
aud[16739]=16'h505;
aud[16740]=16'h4f0;
aud[16741]=16'h4db;
aud[16742]=16'h4c5;
aud[16743]=16'h4b0;
aud[16744]=16'h49b;
aud[16745]=16'h485;
aud[16746]=16'h470;
aud[16747]=16'h45a;
aud[16748]=16'h445;
aud[16749]=16'h430;
aud[16750]=16'h41a;
aud[16751]=16'h405;
aud[16752]=16'h3ef;
aud[16753]=16'h3da;
aud[16754]=16'h3c5;
aud[16755]=16'h3af;
aud[16756]=16'h39a;
aud[16757]=16'h384;
aud[16758]=16'h36f;
aud[16759]=16'h359;
aud[16760]=16'h344;
aud[16761]=16'h32f;
aud[16762]=16'h319;
aud[16763]=16'h304;
aud[16764]=16'h2ee;
aud[16765]=16'h2d9;
aud[16766]=16'h2c4;
aud[16767]=16'h2ae;
aud[16768]=16'h299;
aud[16769]=16'h283;
aud[16770]=16'h26e;
aud[16771]=16'h258;
aud[16772]=16'h243;
aud[16773]=16'h22e;
aud[16774]=16'h218;
aud[16775]=16'h203;
aud[16776]=16'h1ed;
aud[16777]=16'h1d8;
aud[16778]=16'h1c2;
aud[16779]=16'h1ad;
aud[16780]=16'h197;
aud[16781]=16'h182;
aud[16782]=16'h16d;
aud[16783]=16'h157;
aud[16784]=16'h142;
aud[16785]=16'h12c;
aud[16786]=16'h117;
aud[16787]=16'h101;
aud[16788]=16'hec;
aud[16789]=16'hd6;
aud[16790]=16'hc1;
aud[16791]=16'hac;
aud[16792]=16'h96;
aud[16793]=16'h81;
aud[16794]=16'h6b;
aud[16795]=16'h56;
aud[16796]=16'h40;
aud[16797]=16'h2b;
aud[16798]=16'h15;
aud[16799]=16'h0;
aud[16800]=16'hffeb;
aud[16801]=16'hffd5;
aud[16802]=16'hffc0;
aud[16803]=16'hffaa;
aud[16804]=16'hff95;
aud[16805]=16'hff7f;
aud[16806]=16'hff6a;
aud[16807]=16'hff54;
aud[16808]=16'hff3f;
aud[16809]=16'hff2a;
aud[16810]=16'hff14;
aud[16811]=16'hfeff;
aud[16812]=16'hfee9;
aud[16813]=16'hfed4;
aud[16814]=16'hfebe;
aud[16815]=16'hfea9;
aud[16816]=16'hfe93;
aud[16817]=16'hfe7e;
aud[16818]=16'hfe69;
aud[16819]=16'hfe53;
aud[16820]=16'hfe3e;
aud[16821]=16'hfe28;
aud[16822]=16'hfe13;
aud[16823]=16'hfdfd;
aud[16824]=16'hfde8;
aud[16825]=16'hfdd2;
aud[16826]=16'hfdbd;
aud[16827]=16'hfda8;
aud[16828]=16'hfd92;
aud[16829]=16'hfd7d;
aud[16830]=16'hfd67;
aud[16831]=16'hfd52;
aud[16832]=16'hfd3c;
aud[16833]=16'hfd27;
aud[16834]=16'hfd12;
aud[16835]=16'hfcfc;
aud[16836]=16'hfce7;
aud[16837]=16'hfcd1;
aud[16838]=16'hfcbc;
aud[16839]=16'hfca7;
aud[16840]=16'hfc91;
aud[16841]=16'hfc7c;
aud[16842]=16'hfc66;
aud[16843]=16'hfc51;
aud[16844]=16'hfc3b;
aud[16845]=16'hfc26;
aud[16846]=16'hfc11;
aud[16847]=16'hfbfb;
aud[16848]=16'hfbe6;
aud[16849]=16'hfbd0;
aud[16850]=16'hfbbb;
aud[16851]=16'hfba6;
aud[16852]=16'hfb90;
aud[16853]=16'hfb7b;
aud[16854]=16'hfb65;
aud[16855]=16'hfb50;
aud[16856]=16'hfb3b;
aud[16857]=16'hfb25;
aud[16858]=16'hfb10;
aud[16859]=16'hfafb;
aud[16860]=16'hfae5;
aud[16861]=16'hfad0;
aud[16862]=16'hfaba;
aud[16863]=16'hfaa5;
aud[16864]=16'hfa90;
aud[16865]=16'hfa7a;
aud[16866]=16'hfa65;
aud[16867]=16'hfa50;
aud[16868]=16'hfa3a;
aud[16869]=16'hfa25;
aud[16870]=16'hfa0f;
aud[16871]=16'hf9fa;
aud[16872]=16'hf9e5;
aud[16873]=16'hf9cf;
aud[16874]=16'hf9ba;
aud[16875]=16'hf9a5;
aud[16876]=16'hf98f;
aud[16877]=16'hf97a;
aud[16878]=16'hf965;
aud[16879]=16'hf94f;
aud[16880]=16'hf93a;
aud[16881]=16'hf925;
aud[16882]=16'hf90f;
aud[16883]=16'hf8fa;
aud[16884]=16'hf8e5;
aud[16885]=16'hf8cf;
aud[16886]=16'hf8ba;
aud[16887]=16'hf8a5;
aud[16888]=16'hf890;
aud[16889]=16'hf87a;
aud[16890]=16'hf865;
aud[16891]=16'hf850;
aud[16892]=16'hf83a;
aud[16893]=16'hf825;
aud[16894]=16'hf810;
aud[16895]=16'hf7fb;
aud[16896]=16'hf7e5;
aud[16897]=16'hf7d0;
aud[16898]=16'hf7bb;
aud[16899]=16'hf7a5;
aud[16900]=16'hf790;
aud[16901]=16'hf77b;
aud[16902]=16'hf766;
aud[16903]=16'hf750;
aud[16904]=16'hf73b;
aud[16905]=16'hf726;
aud[16906]=16'hf711;
aud[16907]=16'hf6fb;
aud[16908]=16'hf6e6;
aud[16909]=16'hf6d1;
aud[16910]=16'hf6bc;
aud[16911]=16'hf6a7;
aud[16912]=16'hf691;
aud[16913]=16'hf67c;
aud[16914]=16'hf667;
aud[16915]=16'hf652;
aud[16916]=16'hf63d;
aud[16917]=16'hf627;
aud[16918]=16'hf612;
aud[16919]=16'hf5fd;
aud[16920]=16'hf5e8;
aud[16921]=16'hf5d3;
aud[16922]=16'hf5bd;
aud[16923]=16'hf5a8;
aud[16924]=16'hf593;
aud[16925]=16'hf57e;
aud[16926]=16'hf569;
aud[16927]=16'hf554;
aud[16928]=16'hf53f;
aud[16929]=16'hf529;
aud[16930]=16'hf514;
aud[16931]=16'hf4ff;
aud[16932]=16'hf4ea;
aud[16933]=16'hf4d5;
aud[16934]=16'hf4c0;
aud[16935]=16'hf4ab;
aud[16936]=16'hf496;
aud[16937]=16'hf480;
aud[16938]=16'hf46b;
aud[16939]=16'hf456;
aud[16940]=16'hf441;
aud[16941]=16'hf42c;
aud[16942]=16'hf417;
aud[16943]=16'hf402;
aud[16944]=16'hf3ed;
aud[16945]=16'hf3d8;
aud[16946]=16'hf3c3;
aud[16947]=16'hf3ae;
aud[16948]=16'hf399;
aud[16949]=16'hf384;
aud[16950]=16'hf36f;
aud[16951]=16'hf35a;
aud[16952]=16'hf345;
aud[16953]=16'hf330;
aud[16954]=16'hf31b;
aud[16955]=16'hf306;
aud[16956]=16'hf2f1;
aud[16957]=16'hf2dc;
aud[16958]=16'hf2c7;
aud[16959]=16'hf2b2;
aud[16960]=16'hf29d;
aud[16961]=16'hf288;
aud[16962]=16'hf273;
aud[16963]=16'hf25e;
aud[16964]=16'hf249;
aud[16965]=16'hf234;
aud[16966]=16'hf21f;
aud[16967]=16'hf20a;
aud[16968]=16'hf1f5;
aud[16969]=16'hf1e0;
aud[16970]=16'hf1cb;
aud[16971]=16'hf1b6;
aud[16972]=16'hf1a1;
aud[16973]=16'hf18c;
aud[16974]=16'hf178;
aud[16975]=16'hf163;
aud[16976]=16'hf14e;
aud[16977]=16'hf139;
aud[16978]=16'hf124;
aud[16979]=16'hf10f;
aud[16980]=16'hf0fa;
aud[16981]=16'hf0e6;
aud[16982]=16'hf0d1;
aud[16983]=16'hf0bc;
aud[16984]=16'hf0a7;
aud[16985]=16'hf092;
aud[16986]=16'hf07d;
aud[16987]=16'hf069;
aud[16988]=16'hf054;
aud[16989]=16'hf03f;
aud[16990]=16'hf02a;
aud[16991]=16'hf015;
aud[16992]=16'hf001;
aud[16993]=16'hefec;
aud[16994]=16'hefd7;
aud[16995]=16'hefc2;
aud[16996]=16'hefae;
aud[16997]=16'hef99;
aud[16998]=16'hef84;
aud[16999]=16'hef70;
aud[17000]=16'hef5b;
aud[17001]=16'hef46;
aud[17002]=16'hef31;
aud[17003]=16'hef1d;
aud[17004]=16'hef08;
aud[17005]=16'heef3;
aud[17006]=16'heedf;
aud[17007]=16'heeca;
aud[17008]=16'heeb5;
aud[17009]=16'heea1;
aud[17010]=16'hee8c;
aud[17011]=16'hee77;
aud[17012]=16'hee63;
aud[17013]=16'hee4e;
aud[17014]=16'hee3a;
aud[17015]=16'hee25;
aud[17016]=16'hee10;
aud[17017]=16'hedfc;
aud[17018]=16'hede7;
aud[17019]=16'hedd3;
aud[17020]=16'hedbe;
aud[17021]=16'hedaa;
aud[17022]=16'hed95;
aud[17023]=16'hed81;
aud[17024]=16'hed6c;
aud[17025]=16'hed57;
aud[17026]=16'hed43;
aud[17027]=16'hed2e;
aud[17028]=16'hed1a;
aud[17029]=16'hed05;
aud[17030]=16'hecf1;
aud[17031]=16'hecdd;
aud[17032]=16'hecc8;
aud[17033]=16'hecb4;
aud[17034]=16'hec9f;
aud[17035]=16'hec8b;
aud[17036]=16'hec76;
aud[17037]=16'hec62;
aud[17038]=16'hec4d;
aud[17039]=16'hec39;
aud[17040]=16'hec25;
aud[17041]=16'hec10;
aud[17042]=16'hebfc;
aud[17043]=16'hebe8;
aud[17044]=16'hebd3;
aud[17045]=16'hebbf;
aud[17046]=16'hebab;
aud[17047]=16'heb96;
aud[17048]=16'heb82;
aud[17049]=16'heb6e;
aud[17050]=16'heb59;
aud[17051]=16'heb45;
aud[17052]=16'heb31;
aud[17053]=16'heb1c;
aud[17054]=16'heb08;
aud[17055]=16'heaf4;
aud[17056]=16'heae0;
aud[17057]=16'heacb;
aud[17058]=16'heab7;
aud[17059]=16'heaa3;
aud[17060]=16'hea8f;
aud[17061]=16'hea7a;
aud[17062]=16'hea66;
aud[17063]=16'hea52;
aud[17064]=16'hea3e;
aud[17065]=16'hea2a;
aud[17066]=16'hea16;
aud[17067]=16'hea01;
aud[17068]=16'he9ed;
aud[17069]=16'he9d9;
aud[17070]=16'he9c5;
aud[17071]=16'he9b1;
aud[17072]=16'he99d;
aud[17073]=16'he989;
aud[17074]=16'he975;
aud[17075]=16'he961;
aud[17076]=16'he94d;
aud[17077]=16'he939;
aud[17078]=16'he925;
aud[17079]=16'he910;
aud[17080]=16'he8fc;
aud[17081]=16'he8e8;
aud[17082]=16'he8d4;
aud[17083]=16'he8c0;
aud[17084]=16'he8ad;
aud[17085]=16'he899;
aud[17086]=16'he885;
aud[17087]=16'he871;
aud[17088]=16'he85d;
aud[17089]=16'he849;
aud[17090]=16'he835;
aud[17091]=16'he821;
aud[17092]=16'he80d;
aud[17093]=16'he7f9;
aud[17094]=16'he7e5;
aud[17095]=16'he7d1;
aud[17096]=16'he7be;
aud[17097]=16'he7aa;
aud[17098]=16'he796;
aud[17099]=16'he782;
aud[17100]=16'he76e;
aud[17101]=16'he75b;
aud[17102]=16'he747;
aud[17103]=16'he733;
aud[17104]=16'he71f;
aud[17105]=16'he70b;
aud[17106]=16'he6f8;
aud[17107]=16'he6e4;
aud[17108]=16'he6d0;
aud[17109]=16'he6bd;
aud[17110]=16'he6a9;
aud[17111]=16'he695;
aud[17112]=16'he681;
aud[17113]=16'he66e;
aud[17114]=16'he65a;
aud[17115]=16'he646;
aud[17116]=16'he633;
aud[17117]=16'he61f;
aud[17118]=16'he60c;
aud[17119]=16'he5f8;
aud[17120]=16'he5e4;
aud[17121]=16'he5d1;
aud[17122]=16'he5bd;
aud[17123]=16'he5aa;
aud[17124]=16'he596;
aud[17125]=16'he583;
aud[17126]=16'he56f;
aud[17127]=16'he55c;
aud[17128]=16'he548;
aud[17129]=16'he535;
aud[17130]=16'he521;
aud[17131]=16'he50e;
aud[17132]=16'he4fa;
aud[17133]=16'he4e7;
aud[17134]=16'he4d3;
aud[17135]=16'he4c0;
aud[17136]=16'he4ad;
aud[17137]=16'he499;
aud[17138]=16'he486;
aud[17139]=16'he473;
aud[17140]=16'he45f;
aud[17141]=16'he44c;
aud[17142]=16'he438;
aud[17143]=16'he425;
aud[17144]=16'he412;
aud[17145]=16'he3ff;
aud[17146]=16'he3eb;
aud[17147]=16'he3d8;
aud[17148]=16'he3c5;
aud[17149]=16'he3b2;
aud[17150]=16'he39e;
aud[17151]=16'he38b;
aud[17152]=16'he378;
aud[17153]=16'he365;
aud[17154]=16'he352;
aud[17155]=16'he33e;
aud[17156]=16'he32b;
aud[17157]=16'he318;
aud[17158]=16'he305;
aud[17159]=16'he2f2;
aud[17160]=16'he2df;
aud[17161]=16'he2cc;
aud[17162]=16'he2b9;
aud[17163]=16'he2a5;
aud[17164]=16'he292;
aud[17165]=16'he27f;
aud[17166]=16'he26c;
aud[17167]=16'he259;
aud[17168]=16'he246;
aud[17169]=16'he233;
aud[17170]=16'he220;
aud[17171]=16'he20d;
aud[17172]=16'he1fa;
aud[17173]=16'he1e8;
aud[17174]=16'he1d5;
aud[17175]=16'he1c2;
aud[17176]=16'he1af;
aud[17177]=16'he19c;
aud[17178]=16'he189;
aud[17179]=16'he176;
aud[17180]=16'he163;
aud[17181]=16'he151;
aud[17182]=16'he13e;
aud[17183]=16'he12b;
aud[17184]=16'he118;
aud[17185]=16'he105;
aud[17186]=16'he0f3;
aud[17187]=16'he0e0;
aud[17188]=16'he0cd;
aud[17189]=16'he0ba;
aud[17190]=16'he0a8;
aud[17191]=16'he095;
aud[17192]=16'he082;
aud[17193]=16'he070;
aud[17194]=16'he05d;
aud[17195]=16'he04a;
aud[17196]=16'he038;
aud[17197]=16'he025;
aud[17198]=16'he013;
aud[17199]=16'he000;
aud[17200]=16'hdfed;
aud[17201]=16'hdfdb;
aud[17202]=16'hdfc8;
aud[17203]=16'hdfb6;
aud[17204]=16'hdfa3;
aud[17205]=16'hdf91;
aud[17206]=16'hdf7e;
aud[17207]=16'hdf6c;
aud[17208]=16'hdf59;
aud[17209]=16'hdf47;
aud[17210]=16'hdf35;
aud[17211]=16'hdf22;
aud[17212]=16'hdf10;
aud[17213]=16'hdefd;
aud[17214]=16'hdeeb;
aud[17215]=16'hded9;
aud[17216]=16'hdec6;
aud[17217]=16'hdeb4;
aud[17218]=16'hdea2;
aud[17219]=16'hde8f;
aud[17220]=16'hde7d;
aud[17221]=16'hde6b;
aud[17222]=16'hde59;
aud[17223]=16'hde46;
aud[17224]=16'hde34;
aud[17225]=16'hde22;
aud[17226]=16'hde10;
aud[17227]=16'hddfe;
aud[17228]=16'hddeb;
aud[17229]=16'hddd9;
aud[17230]=16'hddc7;
aud[17231]=16'hddb5;
aud[17232]=16'hdda3;
aud[17233]=16'hdd91;
aud[17234]=16'hdd7f;
aud[17235]=16'hdd6d;
aud[17236]=16'hdd5b;
aud[17237]=16'hdd49;
aud[17238]=16'hdd37;
aud[17239]=16'hdd25;
aud[17240]=16'hdd13;
aud[17241]=16'hdd01;
aud[17242]=16'hdcef;
aud[17243]=16'hdcdd;
aud[17244]=16'hdccb;
aud[17245]=16'hdcb9;
aud[17246]=16'hdca7;
aud[17247]=16'hdc95;
aud[17248]=16'hdc83;
aud[17249]=16'hdc72;
aud[17250]=16'hdc60;
aud[17251]=16'hdc4e;
aud[17252]=16'hdc3c;
aud[17253]=16'hdc2a;
aud[17254]=16'hdc19;
aud[17255]=16'hdc07;
aud[17256]=16'hdbf5;
aud[17257]=16'hdbe3;
aud[17258]=16'hdbd2;
aud[17259]=16'hdbc0;
aud[17260]=16'hdbae;
aud[17261]=16'hdb9d;
aud[17262]=16'hdb8b;
aud[17263]=16'hdb79;
aud[17264]=16'hdb68;
aud[17265]=16'hdb56;
aud[17266]=16'hdb45;
aud[17267]=16'hdb33;
aud[17268]=16'hdb22;
aud[17269]=16'hdb10;
aud[17270]=16'hdaff;
aud[17271]=16'hdaed;
aud[17272]=16'hdadc;
aud[17273]=16'hdaca;
aud[17274]=16'hdab9;
aud[17275]=16'hdaa7;
aud[17276]=16'hda96;
aud[17277]=16'hda84;
aud[17278]=16'hda73;
aud[17279]=16'hda62;
aud[17280]=16'hda50;
aud[17281]=16'hda3f;
aud[17282]=16'hda2e;
aud[17283]=16'hda1c;
aud[17284]=16'hda0b;
aud[17285]=16'hd9fa;
aud[17286]=16'hd9e9;
aud[17287]=16'hd9d7;
aud[17288]=16'hd9c6;
aud[17289]=16'hd9b5;
aud[17290]=16'hd9a4;
aud[17291]=16'hd993;
aud[17292]=16'hd982;
aud[17293]=16'hd970;
aud[17294]=16'hd95f;
aud[17295]=16'hd94e;
aud[17296]=16'hd93d;
aud[17297]=16'hd92c;
aud[17298]=16'hd91b;
aud[17299]=16'hd90a;
aud[17300]=16'hd8f9;
aud[17301]=16'hd8e8;
aud[17302]=16'hd8d7;
aud[17303]=16'hd8c6;
aud[17304]=16'hd8b5;
aud[17305]=16'hd8a4;
aud[17306]=16'hd893;
aud[17307]=16'hd882;
aud[17308]=16'hd872;
aud[17309]=16'hd861;
aud[17310]=16'hd850;
aud[17311]=16'hd83f;
aud[17312]=16'hd82e;
aud[17313]=16'hd81e;
aud[17314]=16'hd80d;
aud[17315]=16'hd7fc;
aud[17316]=16'hd7eb;
aud[17317]=16'hd7db;
aud[17318]=16'hd7ca;
aud[17319]=16'hd7b9;
aud[17320]=16'hd7a9;
aud[17321]=16'hd798;
aud[17322]=16'hd787;
aud[17323]=16'hd777;
aud[17324]=16'hd766;
aud[17325]=16'hd756;
aud[17326]=16'hd745;
aud[17327]=16'hd734;
aud[17328]=16'hd724;
aud[17329]=16'hd713;
aud[17330]=16'hd703;
aud[17331]=16'hd6f2;
aud[17332]=16'hd6e2;
aud[17333]=16'hd6d2;
aud[17334]=16'hd6c1;
aud[17335]=16'hd6b1;
aud[17336]=16'hd6a0;
aud[17337]=16'hd690;
aud[17338]=16'hd680;
aud[17339]=16'hd66f;
aud[17340]=16'hd65f;
aud[17341]=16'hd64f;
aud[17342]=16'hd63f;
aud[17343]=16'hd62e;
aud[17344]=16'hd61e;
aud[17345]=16'hd60e;
aud[17346]=16'hd5fe;
aud[17347]=16'hd5ee;
aud[17348]=16'hd5dd;
aud[17349]=16'hd5cd;
aud[17350]=16'hd5bd;
aud[17351]=16'hd5ad;
aud[17352]=16'hd59d;
aud[17353]=16'hd58d;
aud[17354]=16'hd57d;
aud[17355]=16'hd56d;
aud[17356]=16'hd55d;
aud[17357]=16'hd54d;
aud[17358]=16'hd53d;
aud[17359]=16'hd52d;
aud[17360]=16'hd51d;
aud[17361]=16'hd50d;
aud[17362]=16'hd4fd;
aud[17363]=16'hd4ed;
aud[17364]=16'hd4de;
aud[17365]=16'hd4ce;
aud[17366]=16'hd4be;
aud[17367]=16'hd4ae;
aud[17368]=16'hd49e;
aud[17369]=16'hd48f;
aud[17370]=16'hd47f;
aud[17371]=16'hd46f;
aud[17372]=16'hd45f;
aud[17373]=16'hd450;
aud[17374]=16'hd440;
aud[17375]=16'hd430;
aud[17376]=16'hd421;
aud[17377]=16'hd411;
aud[17378]=16'hd402;
aud[17379]=16'hd3f2;
aud[17380]=16'hd3e2;
aud[17381]=16'hd3d3;
aud[17382]=16'hd3c3;
aud[17383]=16'hd3b4;
aud[17384]=16'hd3a4;
aud[17385]=16'hd395;
aud[17386]=16'hd386;
aud[17387]=16'hd376;
aud[17388]=16'hd367;
aud[17389]=16'hd357;
aud[17390]=16'hd348;
aud[17391]=16'hd339;
aud[17392]=16'hd329;
aud[17393]=16'hd31a;
aud[17394]=16'hd30b;
aud[17395]=16'hd2fc;
aud[17396]=16'hd2ec;
aud[17397]=16'hd2dd;
aud[17398]=16'hd2ce;
aud[17399]=16'hd2bf;
aud[17400]=16'hd2b0;
aud[17401]=16'hd2a0;
aud[17402]=16'hd291;
aud[17403]=16'hd282;
aud[17404]=16'hd273;
aud[17405]=16'hd264;
aud[17406]=16'hd255;
aud[17407]=16'hd246;
aud[17408]=16'hd237;
aud[17409]=16'hd228;
aud[17410]=16'hd219;
aud[17411]=16'hd20a;
aud[17412]=16'hd1fb;
aud[17413]=16'hd1ec;
aud[17414]=16'hd1de;
aud[17415]=16'hd1cf;
aud[17416]=16'hd1c0;
aud[17417]=16'hd1b1;
aud[17418]=16'hd1a2;
aud[17419]=16'hd193;
aud[17420]=16'hd185;
aud[17421]=16'hd176;
aud[17422]=16'hd167;
aud[17423]=16'hd159;
aud[17424]=16'hd14a;
aud[17425]=16'hd13b;
aud[17426]=16'hd12d;
aud[17427]=16'hd11e;
aud[17428]=16'hd10f;
aud[17429]=16'hd101;
aud[17430]=16'hd0f2;
aud[17431]=16'hd0e4;
aud[17432]=16'hd0d5;
aud[17433]=16'hd0c7;
aud[17434]=16'hd0b8;
aud[17435]=16'hd0aa;
aud[17436]=16'hd09b;
aud[17437]=16'hd08d;
aud[17438]=16'hd07f;
aud[17439]=16'hd070;
aud[17440]=16'hd062;
aud[17441]=16'hd054;
aud[17442]=16'hd045;
aud[17443]=16'hd037;
aud[17444]=16'hd029;
aud[17445]=16'hd01b;
aud[17446]=16'hd00c;
aud[17447]=16'hcffe;
aud[17448]=16'hcff0;
aud[17449]=16'hcfe2;
aud[17450]=16'hcfd4;
aud[17451]=16'hcfc6;
aud[17452]=16'hcfb8;
aud[17453]=16'hcfa9;
aud[17454]=16'hcf9b;
aud[17455]=16'hcf8d;
aud[17456]=16'hcf7f;
aud[17457]=16'hcf71;
aud[17458]=16'hcf63;
aud[17459]=16'hcf56;
aud[17460]=16'hcf48;
aud[17461]=16'hcf3a;
aud[17462]=16'hcf2c;
aud[17463]=16'hcf1e;
aud[17464]=16'hcf10;
aud[17465]=16'hcf02;
aud[17466]=16'hcef5;
aud[17467]=16'hcee7;
aud[17468]=16'hced9;
aud[17469]=16'hcecb;
aud[17470]=16'hcebe;
aud[17471]=16'hceb0;
aud[17472]=16'hcea2;
aud[17473]=16'hce95;
aud[17474]=16'hce87;
aud[17475]=16'hce79;
aud[17476]=16'hce6c;
aud[17477]=16'hce5e;
aud[17478]=16'hce51;
aud[17479]=16'hce43;
aud[17480]=16'hce36;
aud[17481]=16'hce28;
aud[17482]=16'hce1b;
aud[17483]=16'hce0d;
aud[17484]=16'hce00;
aud[17485]=16'hcdf3;
aud[17486]=16'hcde5;
aud[17487]=16'hcdd8;
aud[17488]=16'hcdcb;
aud[17489]=16'hcdbd;
aud[17490]=16'hcdb0;
aud[17491]=16'hcda3;
aud[17492]=16'hcd96;
aud[17493]=16'hcd88;
aud[17494]=16'hcd7b;
aud[17495]=16'hcd6e;
aud[17496]=16'hcd61;
aud[17497]=16'hcd54;
aud[17498]=16'hcd47;
aud[17499]=16'hcd3a;
aud[17500]=16'hcd2d;
aud[17501]=16'hcd20;
aud[17502]=16'hcd13;
aud[17503]=16'hcd06;
aud[17504]=16'hccf9;
aud[17505]=16'hccec;
aud[17506]=16'hccdf;
aud[17507]=16'hccd2;
aud[17508]=16'hccc5;
aud[17509]=16'hccb8;
aud[17510]=16'hccab;
aud[17511]=16'hcc9f;
aud[17512]=16'hcc92;
aud[17513]=16'hcc85;
aud[17514]=16'hcc78;
aud[17515]=16'hcc6c;
aud[17516]=16'hcc5f;
aud[17517]=16'hcc52;
aud[17518]=16'hcc46;
aud[17519]=16'hcc39;
aud[17520]=16'hcc2c;
aud[17521]=16'hcc20;
aud[17522]=16'hcc13;
aud[17523]=16'hcc07;
aud[17524]=16'hcbfa;
aud[17525]=16'hcbee;
aud[17526]=16'hcbe1;
aud[17527]=16'hcbd5;
aud[17528]=16'hcbc9;
aud[17529]=16'hcbbc;
aud[17530]=16'hcbb0;
aud[17531]=16'hcba3;
aud[17532]=16'hcb97;
aud[17533]=16'hcb8b;
aud[17534]=16'hcb7f;
aud[17535]=16'hcb72;
aud[17536]=16'hcb66;
aud[17537]=16'hcb5a;
aud[17538]=16'hcb4e;
aud[17539]=16'hcb42;
aud[17540]=16'hcb35;
aud[17541]=16'hcb29;
aud[17542]=16'hcb1d;
aud[17543]=16'hcb11;
aud[17544]=16'hcb05;
aud[17545]=16'hcaf9;
aud[17546]=16'hcaed;
aud[17547]=16'hcae1;
aud[17548]=16'hcad5;
aud[17549]=16'hcac9;
aud[17550]=16'hcabd;
aud[17551]=16'hcab1;
aud[17552]=16'hcaa6;
aud[17553]=16'hca9a;
aud[17554]=16'hca8e;
aud[17555]=16'hca82;
aud[17556]=16'hca76;
aud[17557]=16'hca6b;
aud[17558]=16'hca5f;
aud[17559]=16'hca53;
aud[17560]=16'hca48;
aud[17561]=16'hca3c;
aud[17562]=16'hca30;
aud[17563]=16'hca25;
aud[17564]=16'hca19;
aud[17565]=16'hca0e;
aud[17566]=16'hca02;
aud[17567]=16'hc9f7;
aud[17568]=16'hc9eb;
aud[17569]=16'hc9e0;
aud[17570]=16'hc9d4;
aud[17571]=16'hc9c9;
aud[17572]=16'hc9bd;
aud[17573]=16'hc9b2;
aud[17574]=16'hc9a7;
aud[17575]=16'hc99b;
aud[17576]=16'hc990;
aud[17577]=16'hc985;
aud[17578]=16'hc97a;
aud[17579]=16'hc96e;
aud[17580]=16'hc963;
aud[17581]=16'hc958;
aud[17582]=16'hc94d;
aud[17583]=16'hc942;
aud[17584]=16'hc937;
aud[17585]=16'hc92c;
aud[17586]=16'hc920;
aud[17587]=16'hc915;
aud[17588]=16'hc90a;
aud[17589]=16'hc8ff;
aud[17590]=16'hc8f5;
aud[17591]=16'hc8ea;
aud[17592]=16'hc8df;
aud[17593]=16'hc8d4;
aud[17594]=16'hc8c9;
aud[17595]=16'hc8be;
aud[17596]=16'hc8b3;
aud[17597]=16'hc8a9;
aud[17598]=16'hc89e;
aud[17599]=16'hc893;
aud[17600]=16'hc888;
aud[17601]=16'hc87e;
aud[17602]=16'hc873;
aud[17603]=16'hc868;
aud[17604]=16'hc85e;
aud[17605]=16'hc853;
aud[17606]=16'hc849;
aud[17607]=16'hc83e;
aud[17608]=16'hc834;
aud[17609]=16'hc829;
aud[17610]=16'hc81f;
aud[17611]=16'hc814;
aud[17612]=16'hc80a;
aud[17613]=16'hc7ff;
aud[17614]=16'hc7f5;
aud[17615]=16'hc7eb;
aud[17616]=16'hc7e0;
aud[17617]=16'hc7d6;
aud[17618]=16'hc7cc;
aud[17619]=16'hc7c1;
aud[17620]=16'hc7b7;
aud[17621]=16'hc7ad;
aud[17622]=16'hc7a3;
aud[17623]=16'hc799;
aud[17624]=16'hc78f;
aud[17625]=16'hc785;
aud[17626]=16'hc77a;
aud[17627]=16'hc770;
aud[17628]=16'hc766;
aud[17629]=16'hc75c;
aud[17630]=16'hc752;
aud[17631]=16'hc748;
aud[17632]=16'hc73f;
aud[17633]=16'hc735;
aud[17634]=16'hc72b;
aud[17635]=16'hc721;
aud[17636]=16'hc717;
aud[17637]=16'hc70d;
aud[17638]=16'hc703;
aud[17639]=16'hc6fa;
aud[17640]=16'hc6f0;
aud[17641]=16'hc6e6;
aud[17642]=16'hc6dd;
aud[17643]=16'hc6d3;
aud[17644]=16'hc6c9;
aud[17645]=16'hc6c0;
aud[17646]=16'hc6b6;
aud[17647]=16'hc6ad;
aud[17648]=16'hc6a3;
aud[17649]=16'hc69a;
aud[17650]=16'hc690;
aud[17651]=16'hc687;
aud[17652]=16'hc67d;
aud[17653]=16'hc674;
aud[17654]=16'hc66b;
aud[17655]=16'hc661;
aud[17656]=16'hc658;
aud[17657]=16'hc64f;
aud[17658]=16'hc645;
aud[17659]=16'hc63c;
aud[17660]=16'hc633;
aud[17661]=16'hc62a;
aud[17662]=16'hc620;
aud[17663]=16'hc617;
aud[17664]=16'hc60e;
aud[17665]=16'hc605;
aud[17666]=16'hc5fc;
aud[17667]=16'hc5f3;
aud[17668]=16'hc5ea;
aud[17669]=16'hc5e1;
aud[17670]=16'hc5d8;
aud[17671]=16'hc5cf;
aud[17672]=16'hc5c6;
aud[17673]=16'hc5bd;
aud[17674]=16'hc5b4;
aud[17675]=16'hc5ac;
aud[17676]=16'hc5a3;
aud[17677]=16'hc59a;
aud[17678]=16'hc591;
aud[17679]=16'hc588;
aud[17680]=16'hc580;
aud[17681]=16'hc577;
aud[17682]=16'hc56e;
aud[17683]=16'hc566;
aud[17684]=16'hc55d;
aud[17685]=16'hc555;
aud[17686]=16'hc54c;
aud[17687]=16'hc544;
aud[17688]=16'hc53b;
aud[17689]=16'hc533;
aud[17690]=16'hc52a;
aud[17691]=16'hc522;
aud[17692]=16'hc519;
aud[17693]=16'hc511;
aud[17694]=16'hc509;
aud[17695]=16'hc500;
aud[17696]=16'hc4f8;
aud[17697]=16'hc4f0;
aud[17698]=16'hc4e7;
aud[17699]=16'hc4df;
aud[17700]=16'hc4d7;
aud[17701]=16'hc4cf;
aud[17702]=16'hc4c7;
aud[17703]=16'hc4bf;
aud[17704]=16'hc4b6;
aud[17705]=16'hc4ae;
aud[17706]=16'hc4a6;
aud[17707]=16'hc49e;
aud[17708]=16'hc496;
aud[17709]=16'hc48e;
aud[17710]=16'hc486;
aud[17711]=16'hc47f;
aud[17712]=16'hc477;
aud[17713]=16'hc46f;
aud[17714]=16'hc467;
aud[17715]=16'hc45f;
aud[17716]=16'hc457;
aud[17717]=16'hc450;
aud[17718]=16'hc448;
aud[17719]=16'hc440;
aud[17720]=16'hc439;
aud[17721]=16'hc431;
aud[17722]=16'hc429;
aud[17723]=16'hc422;
aud[17724]=16'hc41a;
aud[17725]=16'hc413;
aud[17726]=16'hc40b;
aud[17727]=16'hc404;
aud[17728]=16'hc3fc;
aud[17729]=16'hc3f5;
aud[17730]=16'hc3ed;
aud[17731]=16'hc3e6;
aud[17732]=16'hc3df;
aud[17733]=16'hc3d7;
aud[17734]=16'hc3d0;
aud[17735]=16'hc3c9;
aud[17736]=16'hc3c1;
aud[17737]=16'hc3ba;
aud[17738]=16'hc3b3;
aud[17739]=16'hc3ac;
aud[17740]=16'hc3a5;
aud[17741]=16'hc39d;
aud[17742]=16'hc396;
aud[17743]=16'hc38f;
aud[17744]=16'hc388;
aud[17745]=16'hc381;
aud[17746]=16'hc37a;
aud[17747]=16'hc373;
aud[17748]=16'hc36c;
aud[17749]=16'hc365;
aud[17750]=16'hc35f;
aud[17751]=16'hc358;
aud[17752]=16'hc351;
aud[17753]=16'hc34a;
aud[17754]=16'hc343;
aud[17755]=16'hc33d;
aud[17756]=16'hc336;
aud[17757]=16'hc32f;
aud[17758]=16'hc329;
aud[17759]=16'hc322;
aud[17760]=16'hc31b;
aud[17761]=16'hc315;
aud[17762]=16'hc30e;
aud[17763]=16'hc308;
aud[17764]=16'hc301;
aud[17765]=16'hc2fb;
aud[17766]=16'hc2f4;
aud[17767]=16'hc2ee;
aud[17768]=16'hc2e7;
aud[17769]=16'hc2e1;
aud[17770]=16'hc2db;
aud[17771]=16'hc2d4;
aud[17772]=16'hc2ce;
aud[17773]=16'hc2c8;
aud[17774]=16'hc2c1;
aud[17775]=16'hc2bb;
aud[17776]=16'hc2b5;
aud[17777]=16'hc2af;
aud[17778]=16'hc2a9;
aud[17779]=16'hc2a3;
aud[17780]=16'hc29d;
aud[17781]=16'hc297;
aud[17782]=16'hc291;
aud[17783]=16'hc28b;
aud[17784]=16'hc285;
aud[17785]=16'hc27f;
aud[17786]=16'hc279;
aud[17787]=16'hc273;
aud[17788]=16'hc26d;
aud[17789]=16'hc267;
aud[17790]=16'hc261;
aud[17791]=16'hc25c;
aud[17792]=16'hc256;
aud[17793]=16'hc250;
aud[17794]=16'hc24a;
aud[17795]=16'hc245;
aud[17796]=16'hc23f;
aud[17797]=16'hc239;
aud[17798]=16'hc234;
aud[17799]=16'hc22e;
aud[17800]=16'hc229;
aud[17801]=16'hc223;
aud[17802]=16'hc21e;
aud[17803]=16'hc218;
aud[17804]=16'hc213;
aud[17805]=16'hc20d;
aud[17806]=16'hc208;
aud[17807]=16'hc203;
aud[17808]=16'hc1fd;
aud[17809]=16'hc1f8;
aud[17810]=16'hc1f3;
aud[17811]=16'hc1ee;
aud[17812]=16'hc1e8;
aud[17813]=16'hc1e3;
aud[17814]=16'hc1de;
aud[17815]=16'hc1d9;
aud[17816]=16'hc1d4;
aud[17817]=16'hc1cf;
aud[17818]=16'hc1ca;
aud[17819]=16'hc1c5;
aud[17820]=16'hc1c0;
aud[17821]=16'hc1bb;
aud[17822]=16'hc1b6;
aud[17823]=16'hc1b1;
aud[17824]=16'hc1ac;
aud[17825]=16'hc1a7;
aud[17826]=16'hc1a2;
aud[17827]=16'hc19e;
aud[17828]=16'hc199;
aud[17829]=16'hc194;
aud[17830]=16'hc18f;
aud[17831]=16'hc18b;
aud[17832]=16'hc186;
aud[17833]=16'hc181;
aud[17834]=16'hc17d;
aud[17835]=16'hc178;
aud[17836]=16'hc174;
aud[17837]=16'hc16f;
aud[17838]=16'hc16b;
aud[17839]=16'hc166;
aud[17840]=16'hc162;
aud[17841]=16'hc15d;
aud[17842]=16'hc159;
aud[17843]=16'hc154;
aud[17844]=16'hc150;
aud[17845]=16'hc14c;
aud[17846]=16'hc147;
aud[17847]=16'hc143;
aud[17848]=16'hc13f;
aud[17849]=16'hc13b;
aud[17850]=16'hc137;
aud[17851]=16'hc133;
aud[17852]=16'hc12e;
aud[17853]=16'hc12a;
aud[17854]=16'hc126;
aud[17855]=16'hc122;
aud[17856]=16'hc11e;
aud[17857]=16'hc11a;
aud[17858]=16'hc116;
aud[17859]=16'hc112;
aud[17860]=16'hc10e;
aud[17861]=16'hc10b;
aud[17862]=16'hc107;
aud[17863]=16'hc103;
aud[17864]=16'hc0ff;
aud[17865]=16'hc0fb;
aud[17866]=16'hc0f8;
aud[17867]=16'hc0f4;
aud[17868]=16'hc0f0;
aud[17869]=16'hc0ed;
aud[17870]=16'hc0e9;
aud[17871]=16'hc0e5;
aud[17872]=16'hc0e2;
aud[17873]=16'hc0de;
aud[17874]=16'hc0db;
aud[17875]=16'hc0d7;
aud[17876]=16'hc0d4;
aud[17877]=16'hc0d0;
aud[17878]=16'hc0cd;
aud[17879]=16'hc0ca;
aud[17880]=16'hc0c6;
aud[17881]=16'hc0c3;
aud[17882]=16'hc0c0;
aud[17883]=16'hc0bd;
aud[17884]=16'hc0b9;
aud[17885]=16'hc0b6;
aud[17886]=16'hc0b3;
aud[17887]=16'hc0b0;
aud[17888]=16'hc0ad;
aud[17889]=16'hc0aa;
aud[17890]=16'hc0a6;
aud[17891]=16'hc0a3;
aud[17892]=16'hc0a0;
aud[17893]=16'hc09d;
aud[17894]=16'hc09b;
aud[17895]=16'hc098;
aud[17896]=16'hc095;
aud[17897]=16'hc092;
aud[17898]=16'hc08f;
aud[17899]=16'hc08c;
aud[17900]=16'hc089;
aud[17901]=16'hc087;
aud[17902]=16'hc084;
aud[17903]=16'hc081;
aud[17904]=16'hc07f;
aud[17905]=16'hc07c;
aud[17906]=16'hc079;
aud[17907]=16'hc077;
aud[17908]=16'hc074;
aud[17909]=16'hc072;
aud[17910]=16'hc06f;
aud[17911]=16'hc06d;
aud[17912]=16'hc06a;
aud[17913]=16'hc068;
aud[17914]=16'hc065;
aud[17915]=16'hc063;
aud[17916]=16'hc061;
aud[17917]=16'hc05e;
aud[17918]=16'hc05c;
aud[17919]=16'hc05a;
aud[17920]=16'hc058;
aud[17921]=16'hc055;
aud[17922]=16'hc053;
aud[17923]=16'hc051;
aud[17924]=16'hc04f;
aud[17925]=16'hc04d;
aud[17926]=16'hc04b;
aud[17927]=16'hc049;
aud[17928]=16'hc047;
aud[17929]=16'hc045;
aud[17930]=16'hc043;
aud[17931]=16'hc041;
aud[17932]=16'hc03f;
aud[17933]=16'hc03d;
aud[17934]=16'hc03b;
aud[17935]=16'hc039;
aud[17936]=16'hc038;
aud[17937]=16'hc036;
aud[17938]=16'hc034;
aud[17939]=16'hc033;
aud[17940]=16'hc031;
aud[17941]=16'hc02f;
aud[17942]=16'hc02e;
aud[17943]=16'hc02c;
aud[17944]=16'hc02a;
aud[17945]=16'hc029;
aud[17946]=16'hc027;
aud[17947]=16'hc026;
aud[17948]=16'hc024;
aud[17949]=16'hc023;
aud[17950]=16'hc022;
aud[17951]=16'hc020;
aud[17952]=16'hc01f;
aud[17953]=16'hc01e;
aud[17954]=16'hc01c;
aud[17955]=16'hc01b;
aud[17956]=16'hc01a;
aud[17957]=16'hc019;
aud[17958]=16'hc018;
aud[17959]=16'hc016;
aud[17960]=16'hc015;
aud[17961]=16'hc014;
aud[17962]=16'hc013;
aud[17963]=16'hc012;
aud[17964]=16'hc011;
aud[17965]=16'hc010;
aud[17966]=16'hc00f;
aud[17967]=16'hc00e;
aud[17968]=16'hc00d;
aud[17969]=16'hc00d;
aud[17970]=16'hc00c;
aud[17971]=16'hc00b;
aud[17972]=16'hc00a;
aud[17973]=16'hc009;
aud[17974]=16'hc009;
aud[17975]=16'hc008;
aud[17976]=16'hc007;
aud[17977]=16'hc007;
aud[17978]=16'hc006;
aud[17979]=16'hc006;
aud[17980]=16'hc005;
aud[17981]=16'hc005;
aud[17982]=16'hc004;
aud[17983]=16'hc004;
aud[17984]=16'hc003;
aud[17985]=16'hc003;
aud[17986]=16'hc002;
aud[17987]=16'hc002;
aud[17988]=16'hc002;
aud[17989]=16'hc001;
aud[17990]=16'hc001;
aud[17991]=16'hc001;
aud[17992]=16'hc001;
aud[17993]=16'hc001;
aud[17994]=16'hc000;
aud[17995]=16'hc000;
aud[17996]=16'hc000;
aud[17997]=16'hc000;
aud[17998]=16'hc000;
aud[17999]=16'hc000;
aud[18000]=16'hc000;
aud[18001]=16'hc000;
aud[18002]=16'hc000;
aud[18003]=16'hc000;
aud[18004]=16'hc000;
aud[18005]=16'hc001;
aud[18006]=16'hc001;
aud[18007]=16'hc001;
aud[18008]=16'hc001;
aud[18009]=16'hc001;
aud[18010]=16'hc002;
aud[18011]=16'hc002;
aud[18012]=16'hc002;
aud[18013]=16'hc003;
aud[18014]=16'hc003;
aud[18015]=16'hc004;
aud[18016]=16'hc004;
aud[18017]=16'hc005;
aud[18018]=16'hc005;
aud[18019]=16'hc006;
aud[18020]=16'hc006;
aud[18021]=16'hc007;
aud[18022]=16'hc007;
aud[18023]=16'hc008;
aud[18024]=16'hc009;
aud[18025]=16'hc009;
aud[18026]=16'hc00a;
aud[18027]=16'hc00b;
aud[18028]=16'hc00c;
aud[18029]=16'hc00d;
aud[18030]=16'hc00d;
aud[18031]=16'hc00e;
aud[18032]=16'hc00f;
aud[18033]=16'hc010;
aud[18034]=16'hc011;
aud[18035]=16'hc012;
aud[18036]=16'hc013;
aud[18037]=16'hc014;
aud[18038]=16'hc015;
aud[18039]=16'hc016;
aud[18040]=16'hc018;
aud[18041]=16'hc019;
aud[18042]=16'hc01a;
aud[18043]=16'hc01b;
aud[18044]=16'hc01c;
aud[18045]=16'hc01e;
aud[18046]=16'hc01f;
aud[18047]=16'hc020;
aud[18048]=16'hc022;
aud[18049]=16'hc023;
aud[18050]=16'hc024;
aud[18051]=16'hc026;
aud[18052]=16'hc027;
aud[18053]=16'hc029;
aud[18054]=16'hc02a;
aud[18055]=16'hc02c;
aud[18056]=16'hc02e;
aud[18057]=16'hc02f;
aud[18058]=16'hc031;
aud[18059]=16'hc033;
aud[18060]=16'hc034;
aud[18061]=16'hc036;
aud[18062]=16'hc038;
aud[18063]=16'hc039;
aud[18064]=16'hc03b;
aud[18065]=16'hc03d;
aud[18066]=16'hc03f;
aud[18067]=16'hc041;
aud[18068]=16'hc043;
aud[18069]=16'hc045;
aud[18070]=16'hc047;
aud[18071]=16'hc049;
aud[18072]=16'hc04b;
aud[18073]=16'hc04d;
aud[18074]=16'hc04f;
aud[18075]=16'hc051;
aud[18076]=16'hc053;
aud[18077]=16'hc055;
aud[18078]=16'hc058;
aud[18079]=16'hc05a;
aud[18080]=16'hc05c;
aud[18081]=16'hc05e;
aud[18082]=16'hc061;
aud[18083]=16'hc063;
aud[18084]=16'hc065;
aud[18085]=16'hc068;
aud[18086]=16'hc06a;
aud[18087]=16'hc06d;
aud[18088]=16'hc06f;
aud[18089]=16'hc072;
aud[18090]=16'hc074;
aud[18091]=16'hc077;
aud[18092]=16'hc079;
aud[18093]=16'hc07c;
aud[18094]=16'hc07f;
aud[18095]=16'hc081;
aud[18096]=16'hc084;
aud[18097]=16'hc087;
aud[18098]=16'hc089;
aud[18099]=16'hc08c;
aud[18100]=16'hc08f;
aud[18101]=16'hc092;
aud[18102]=16'hc095;
aud[18103]=16'hc098;
aud[18104]=16'hc09b;
aud[18105]=16'hc09d;
aud[18106]=16'hc0a0;
aud[18107]=16'hc0a3;
aud[18108]=16'hc0a6;
aud[18109]=16'hc0aa;
aud[18110]=16'hc0ad;
aud[18111]=16'hc0b0;
aud[18112]=16'hc0b3;
aud[18113]=16'hc0b6;
aud[18114]=16'hc0b9;
aud[18115]=16'hc0bd;
aud[18116]=16'hc0c0;
aud[18117]=16'hc0c3;
aud[18118]=16'hc0c6;
aud[18119]=16'hc0ca;
aud[18120]=16'hc0cd;
aud[18121]=16'hc0d0;
aud[18122]=16'hc0d4;
aud[18123]=16'hc0d7;
aud[18124]=16'hc0db;
aud[18125]=16'hc0de;
aud[18126]=16'hc0e2;
aud[18127]=16'hc0e5;
aud[18128]=16'hc0e9;
aud[18129]=16'hc0ed;
aud[18130]=16'hc0f0;
aud[18131]=16'hc0f4;
aud[18132]=16'hc0f8;
aud[18133]=16'hc0fb;
aud[18134]=16'hc0ff;
aud[18135]=16'hc103;
aud[18136]=16'hc107;
aud[18137]=16'hc10b;
aud[18138]=16'hc10e;
aud[18139]=16'hc112;
aud[18140]=16'hc116;
aud[18141]=16'hc11a;
aud[18142]=16'hc11e;
aud[18143]=16'hc122;
aud[18144]=16'hc126;
aud[18145]=16'hc12a;
aud[18146]=16'hc12e;
aud[18147]=16'hc133;
aud[18148]=16'hc137;
aud[18149]=16'hc13b;
aud[18150]=16'hc13f;
aud[18151]=16'hc143;
aud[18152]=16'hc147;
aud[18153]=16'hc14c;
aud[18154]=16'hc150;
aud[18155]=16'hc154;
aud[18156]=16'hc159;
aud[18157]=16'hc15d;
aud[18158]=16'hc162;
aud[18159]=16'hc166;
aud[18160]=16'hc16b;
aud[18161]=16'hc16f;
aud[18162]=16'hc174;
aud[18163]=16'hc178;
aud[18164]=16'hc17d;
aud[18165]=16'hc181;
aud[18166]=16'hc186;
aud[18167]=16'hc18b;
aud[18168]=16'hc18f;
aud[18169]=16'hc194;
aud[18170]=16'hc199;
aud[18171]=16'hc19e;
aud[18172]=16'hc1a2;
aud[18173]=16'hc1a7;
aud[18174]=16'hc1ac;
aud[18175]=16'hc1b1;
aud[18176]=16'hc1b6;
aud[18177]=16'hc1bb;
aud[18178]=16'hc1c0;
aud[18179]=16'hc1c5;
aud[18180]=16'hc1ca;
aud[18181]=16'hc1cf;
aud[18182]=16'hc1d4;
aud[18183]=16'hc1d9;
aud[18184]=16'hc1de;
aud[18185]=16'hc1e3;
aud[18186]=16'hc1e8;
aud[18187]=16'hc1ee;
aud[18188]=16'hc1f3;
aud[18189]=16'hc1f8;
aud[18190]=16'hc1fd;
aud[18191]=16'hc203;
aud[18192]=16'hc208;
aud[18193]=16'hc20d;
aud[18194]=16'hc213;
aud[18195]=16'hc218;
aud[18196]=16'hc21e;
aud[18197]=16'hc223;
aud[18198]=16'hc229;
aud[18199]=16'hc22e;
aud[18200]=16'hc234;
aud[18201]=16'hc239;
aud[18202]=16'hc23f;
aud[18203]=16'hc245;
aud[18204]=16'hc24a;
aud[18205]=16'hc250;
aud[18206]=16'hc256;
aud[18207]=16'hc25c;
aud[18208]=16'hc261;
aud[18209]=16'hc267;
aud[18210]=16'hc26d;
aud[18211]=16'hc273;
aud[18212]=16'hc279;
aud[18213]=16'hc27f;
aud[18214]=16'hc285;
aud[18215]=16'hc28b;
aud[18216]=16'hc291;
aud[18217]=16'hc297;
aud[18218]=16'hc29d;
aud[18219]=16'hc2a3;
aud[18220]=16'hc2a9;
aud[18221]=16'hc2af;
aud[18222]=16'hc2b5;
aud[18223]=16'hc2bb;
aud[18224]=16'hc2c1;
aud[18225]=16'hc2c8;
aud[18226]=16'hc2ce;
aud[18227]=16'hc2d4;
aud[18228]=16'hc2db;
aud[18229]=16'hc2e1;
aud[18230]=16'hc2e7;
aud[18231]=16'hc2ee;
aud[18232]=16'hc2f4;
aud[18233]=16'hc2fb;
aud[18234]=16'hc301;
aud[18235]=16'hc308;
aud[18236]=16'hc30e;
aud[18237]=16'hc315;
aud[18238]=16'hc31b;
aud[18239]=16'hc322;
aud[18240]=16'hc329;
aud[18241]=16'hc32f;
aud[18242]=16'hc336;
aud[18243]=16'hc33d;
aud[18244]=16'hc343;
aud[18245]=16'hc34a;
aud[18246]=16'hc351;
aud[18247]=16'hc358;
aud[18248]=16'hc35f;
aud[18249]=16'hc365;
aud[18250]=16'hc36c;
aud[18251]=16'hc373;
aud[18252]=16'hc37a;
aud[18253]=16'hc381;
aud[18254]=16'hc388;
aud[18255]=16'hc38f;
aud[18256]=16'hc396;
aud[18257]=16'hc39d;
aud[18258]=16'hc3a5;
aud[18259]=16'hc3ac;
aud[18260]=16'hc3b3;
aud[18261]=16'hc3ba;
aud[18262]=16'hc3c1;
aud[18263]=16'hc3c9;
aud[18264]=16'hc3d0;
aud[18265]=16'hc3d7;
aud[18266]=16'hc3df;
aud[18267]=16'hc3e6;
aud[18268]=16'hc3ed;
aud[18269]=16'hc3f5;
aud[18270]=16'hc3fc;
aud[18271]=16'hc404;
aud[18272]=16'hc40b;
aud[18273]=16'hc413;
aud[18274]=16'hc41a;
aud[18275]=16'hc422;
aud[18276]=16'hc429;
aud[18277]=16'hc431;
aud[18278]=16'hc439;
aud[18279]=16'hc440;
aud[18280]=16'hc448;
aud[18281]=16'hc450;
aud[18282]=16'hc457;
aud[18283]=16'hc45f;
aud[18284]=16'hc467;
aud[18285]=16'hc46f;
aud[18286]=16'hc477;
aud[18287]=16'hc47f;
aud[18288]=16'hc486;
aud[18289]=16'hc48e;
aud[18290]=16'hc496;
aud[18291]=16'hc49e;
aud[18292]=16'hc4a6;
aud[18293]=16'hc4ae;
aud[18294]=16'hc4b6;
aud[18295]=16'hc4bf;
aud[18296]=16'hc4c7;
aud[18297]=16'hc4cf;
aud[18298]=16'hc4d7;
aud[18299]=16'hc4df;
aud[18300]=16'hc4e7;
aud[18301]=16'hc4f0;
aud[18302]=16'hc4f8;
aud[18303]=16'hc500;
aud[18304]=16'hc509;
aud[18305]=16'hc511;
aud[18306]=16'hc519;
aud[18307]=16'hc522;
aud[18308]=16'hc52a;
aud[18309]=16'hc533;
aud[18310]=16'hc53b;
aud[18311]=16'hc544;
aud[18312]=16'hc54c;
aud[18313]=16'hc555;
aud[18314]=16'hc55d;
aud[18315]=16'hc566;
aud[18316]=16'hc56e;
aud[18317]=16'hc577;
aud[18318]=16'hc580;
aud[18319]=16'hc588;
aud[18320]=16'hc591;
aud[18321]=16'hc59a;
aud[18322]=16'hc5a3;
aud[18323]=16'hc5ac;
aud[18324]=16'hc5b4;
aud[18325]=16'hc5bd;
aud[18326]=16'hc5c6;
aud[18327]=16'hc5cf;
aud[18328]=16'hc5d8;
aud[18329]=16'hc5e1;
aud[18330]=16'hc5ea;
aud[18331]=16'hc5f3;
aud[18332]=16'hc5fc;
aud[18333]=16'hc605;
aud[18334]=16'hc60e;
aud[18335]=16'hc617;
aud[18336]=16'hc620;
aud[18337]=16'hc62a;
aud[18338]=16'hc633;
aud[18339]=16'hc63c;
aud[18340]=16'hc645;
aud[18341]=16'hc64f;
aud[18342]=16'hc658;
aud[18343]=16'hc661;
aud[18344]=16'hc66b;
aud[18345]=16'hc674;
aud[18346]=16'hc67d;
aud[18347]=16'hc687;
aud[18348]=16'hc690;
aud[18349]=16'hc69a;
aud[18350]=16'hc6a3;
aud[18351]=16'hc6ad;
aud[18352]=16'hc6b6;
aud[18353]=16'hc6c0;
aud[18354]=16'hc6c9;
aud[18355]=16'hc6d3;
aud[18356]=16'hc6dd;
aud[18357]=16'hc6e6;
aud[18358]=16'hc6f0;
aud[18359]=16'hc6fa;
aud[18360]=16'hc703;
aud[18361]=16'hc70d;
aud[18362]=16'hc717;
aud[18363]=16'hc721;
aud[18364]=16'hc72b;
aud[18365]=16'hc735;
aud[18366]=16'hc73f;
aud[18367]=16'hc748;
aud[18368]=16'hc752;
aud[18369]=16'hc75c;
aud[18370]=16'hc766;
aud[18371]=16'hc770;
aud[18372]=16'hc77a;
aud[18373]=16'hc785;
aud[18374]=16'hc78f;
aud[18375]=16'hc799;
aud[18376]=16'hc7a3;
aud[18377]=16'hc7ad;
aud[18378]=16'hc7b7;
aud[18379]=16'hc7c1;
aud[18380]=16'hc7cc;
aud[18381]=16'hc7d6;
aud[18382]=16'hc7e0;
aud[18383]=16'hc7eb;
aud[18384]=16'hc7f5;
aud[18385]=16'hc7ff;
aud[18386]=16'hc80a;
aud[18387]=16'hc814;
aud[18388]=16'hc81f;
aud[18389]=16'hc829;
aud[18390]=16'hc834;
aud[18391]=16'hc83e;
aud[18392]=16'hc849;
aud[18393]=16'hc853;
aud[18394]=16'hc85e;
aud[18395]=16'hc868;
aud[18396]=16'hc873;
aud[18397]=16'hc87e;
aud[18398]=16'hc888;
aud[18399]=16'hc893;
aud[18400]=16'hc89e;
aud[18401]=16'hc8a9;
aud[18402]=16'hc8b3;
aud[18403]=16'hc8be;
aud[18404]=16'hc8c9;
aud[18405]=16'hc8d4;
aud[18406]=16'hc8df;
aud[18407]=16'hc8ea;
aud[18408]=16'hc8f5;
aud[18409]=16'hc8ff;
aud[18410]=16'hc90a;
aud[18411]=16'hc915;
aud[18412]=16'hc920;
aud[18413]=16'hc92c;
aud[18414]=16'hc937;
aud[18415]=16'hc942;
aud[18416]=16'hc94d;
aud[18417]=16'hc958;
aud[18418]=16'hc963;
aud[18419]=16'hc96e;
aud[18420]=16'hc97a;
aud[18421]=16'hc985;
aud[18422]=16'hc990;
aud[18423]=16'hc99b;
aud[18424]=16'hc9a7;
aud[18425]=16'hc9b2;
aud[18426]=16'hc9bd;
aud[18427]=16'hc9c9;
aud[18428]=16'hc9d4;
aud[18429]=16'hc9e0;
aud[18430]=16'hc9eb;
aud[18431]=16'hc9f7;
aud[18432]=16'hca02;
aud[18433]=16'hca0e;
aud[18434]=16'hca19;
aud[18435]=16'hca25;
aud[18436]=16'hca30;
aud[18437]=16'hca3c;
aud[18438]=16'hca48;
aud[18439]=16'hca53;
aud[18440]=16'hca5f;
aud[18441]=16'hca6b;
aud[18442]=16'hca76;
aud[18443]=16'hca82;
aud[18444]=16'hca8e;
aud[18445]=16'hca9a;
aud[18446]=16'hcaa6;
aud[18447]=16'hcab1;
aud[18448]=16'hcabd;
aud[18449]=16'hcac9;
aud[18450]=16'hcad5;
aud[18451]=16'hcae1;
aud[18452]=16'hcaed;
aud[18453]=16'hcaf9;
aud[18454]=16'hcb05;
aud[18455]=16'hcb11;
aud[18456]=16'hcb1d;
aud[18457]=16'hcb29;
aud[18458]=16'hcb35;
aud[18459]=16'hcb42;
aud[18460]=16'hcb4e;
aud[18461]=16'hcb5a;
aud[18462]=16'hcb66;
aud[18463]=16'hcb72;
aud[18464]=16'hcb7f;
aud[18465]=16'hcb8b;
aud[18466]=16'hcb97;
aud[18467]=16'hcba3;
aud[18468]=16'hcbb0;
aud[18469]=16'hcbbc;
aud[18470]=16'hcbc9;
aud[18471]=16'hcbd5;
aud[18472]=16'hcbe1;
aud[18473]=16'hcbee;
aud[18474]=16'hcbfa;
aud[18475]=16'hcc07;
aud[18476]=16'hcc13;
aud[18477]=16'hcc20;
aud[18478]=16'hcc2c;
aud[18479]=16'hcc39;
aud[18480]=16'hcc46;
aud[18481]=16'hcc52;
aud[18482]=16'hcc5f;
aud[18483]=16'hcc6c;
aud[18484]=16'hcc78;
aud[18485]=16'hcc85;
aud[18486]=16'hcc92;
aud[18487]=16'hcc9f;
aud[18488]=16'hccab;
aud[18489]=16'hccb8;
aud[18490]=16'hccc5;
aud[18491]=16'hccd2;
aud[18492]=16'hccdf;
aud[18493]=16'hccec;
aud[18494]=16'hccf9;
aud[18495]=16'hcd06;
aud[18496]=16'hcd13;
aud[18497]=16'hcd20;
aud[18498]=16'hcd2d;
aud[18499]=16'hcd3a;
aud[18500]=16'hcd47;
aud[18501]=16'hcd54;
aud[18502]=16'hcd61;
aud[18503]=16'hcd6e;
aud[18504]=16'hcd7b;
aud[18505]=16'hcd88;
aud[18506]=16'hcd96;
aud[18507]=16'hcda3;
aud[18508]=16'hcdb0;
aud[18509]=16'hcdbd;
aud[18510]=16'hcdcb;
aud[18511]=16'hcdd8;
aud[18512]=16'hcde5;
aud[18513]=16'hcdf3;
aud[18514]=16'hce00;
aud[18515]=16'hce0d;
aud[18516]=16'hce1b;
aud[18517]=16'hce28;
aud[18518]=16'hce36;
aud[18519]=16'hce43;
aud[18520]=16'hce51;
aud[18521]=16'hce5e;
aud[18522]=16'hce6c;
aud[18523]=16'hce79;
aud[18524]=16'hce87;
aud[18525]=16'hce95;
aud[18526]=16'hcea2;
aud[18527]=16'hceb0;
aud[18528]=16'hcebe;
aud[18529]=16'hcecb;
aud[18530]=16'hced9;
aud[18531]=16'hcee7;
aud[18532]=16'hcef5;
aud[18533]=16'hcf02;
aud[18534]=16'hcf10;
aud[18535]=16'hcf1e;
aud[18536]=16'hcf2c;
aud[18537]=16'hcf3a;
aud[18538]=16'hcf48;
aud[18539]=16'hcf56;
aud[18540]=16'hcf63;
aud[18541]=16'hcf71;
aud[18542]=16'hcf7f;
aud[18543]=16'hcf8d;
aud[18544]=16'hcf9b;
aud[18545]=16'hcfa9;
aud[18546]=16'hcfb8;
aud[18547]=16'hcfc6;
aud[18548]=16'hcfd4;
aud[18549]=16'hcfe2;
aud[18550]=16'hcff0;
aud[18551]=16'hcffe;
aud[18552]=16'hd00c;
aud[18553]=16'hd01b;
aud[18554]=16'hd029;
aud[18555]=16'hd037;
aud[18556]=16'hd045;
aud[18557]=16'hd054;
aud[18558]=16'hd062;
aud[18559]=16'hd070;
aud[18560]=16'hd07f;
aud[18561]=16'hd08d;
aud[18562]=16'hd09b;
aud[18563]=16'hd0aa;
aud[18564]=16'hd0b8;
aud[18565]=16'hd0c7;
aud[18566]=16'hd0d5;
aud[18567]=16'hd0e4;
aud[18568]=16'hd0f2;
aud[18569]=16'hd101;
aud[18570]=16'hd10f;
aud[18571]=16'hd11e;
aud[18572]=16'hd12d;
aud[18573]=16'hd13b;
aud[18574]=16'hd14a;
aud[18575]=16'hd159;
aud[18576]=16'hd167;
aud[18577]=16'hd176;
aud[18578]=16'hd185;
aud[18579]=16'hd193;
aud[18580]=16'hd1a2;
aud[18581]=16'hd1b1;
aud[18582]=16'hd1c0;
aud[18583]=16'hd1cf;
aud[18584]=16'hd1de;
aud[18585]=16'hd1ec;
aud[18586]=16'hd1fb;
aud[18587]=16'hd20a;
aud[18588]=16'hd219;
aud[18589]=16'hd228;
aud[18590]=16'hd237;
aud[18591]=16'hd246;
aud[18592]=16'hd255;
aud[18593]=16'hd264;
aud[18594]=16'hd273;
aud[18595]=16'hd282;
aud[18596]=16'hd291;
aud[18597]=16'hd2a0;
aud[18598]=16'hd2b0;
aud[18599]=16'hd2bf;
aud[18600]=16'hd2ce;
aud[18601]=16'hd2dd;
aud[18602]=16'hd2ec;
aud[18603]=16'hd2fc;
aud[18604]=16'hd30b;
aud[18605]=16'hd31a;
aud[18606]=16'hd329;
aud[18607]=16'hd339;
aud[18608]=16'hd348;
aud[18609]=16'hd357;
aud[18610]=16'hd367;
aud[18611]=16'hd376;
aud[18612]=16'hd386;
aud[18613]=16'hd395;
aud[18614]=16'hd3a4;
aud[18615]=16'hd3b4;
aud[18616]=16'hd3c3;
aud[18617]=16'hd3d3;
aud[18618]=16'hd3e2;
aud[18619]=16'hd3f2;
aud[18620]=16'hd402;
aud[18621]=16'hd411;
aud[18622]=16'hd421;
aud[18623]=16'hd430;
aud[18624]=16'hd440;
aud[18625]=16'hd450;
aud[18626]=16'hd45f;
aud[18627]=16'hd46f;
aud[18628]=16'hd47f;
aud[18629]=16'hd48f;
aud[18630]=16'hd49e;
aud[18631]=16'hd4ae;
aud[18632]=16'hd4be;
aud[18633]=16'hd4ce;
aud[18634]=16'hd4de;
aud[18635]=16'hd4ed;
aud[18636]=16'hd4fd;
aud[18637]=16'hd50d;
aud[18638]=16'hd51d;
aud[18639]=16'hd52d;
aud[18640]=16'hd53d;
aud[18641]=16'hd54d;
aud[18642]=16'hd55d;
aud[18643]=16'hd56d;
aud[18644]=16'hd57d;
aud[18645]=16'hd58d;
aud[18646]=16'hd59d;
aud[18647]=16'hd5ad;
aud[18648]=16'hd5bd;
aud[18649]=16'hd5cd;
aud[18650]=16'hd5dd;
aud[18651]=16'hd5ee;
aud[18652]=16'hd5fe;
aud[18653]=16'hd60e;
aud[18654]=16'hd61e;
aud[18655]=16'hd62e;
aud[18656]=16'hd63f;
aud[18657]=16'hd64f;
aud[18658]=16'hd65f;
aud[18659]=16'hd66f;
aud[18660]=16'hd680;
aud[18661]=16'hd690;
aud[18662]=16'hd6a0;
aud[18663]=16'hd6b1;
aud[18664]=16'hd6c1;
aud[18665]=16'hd6d2;
aud[18666]=16'hd6e2;
aud[18667]=16'hd6f2;
aud[18668]=16'hd703;
aud[18669]=16'hd713;
aud[18670]=16'hd724;
aud[18671]=16'hd734;
aud[18672]=16'hd745;
aud[18673]=16'hd756;
aud[18674]=16'hd766;
aud[18675]=16'hd777;
aud[18676]=16'hd787;
aud[18677]=16'hd798;
aud[18678]=16'hd7a9;
aud[18679]=16'hd7b9;
aud[18680]=16'hd7ca;
aud[18681]=16'hd7db;
aud[18682]=16'hd7eb;
aud[18683]=16'hd7fc;
aud[18684]=16'hd80d;
aud[18685]=16'hd81e;
aud[18686]=16'hd82e;
aud[18687]=16'hd83f;
aud[18688]=16'hd850;
aud[18689]=16'hd861;
aud[18690]=16'hd872;
aud[18691]=16'hd882;
aud[18692]=16'hd893;
aud[18693]=16'hd8a4;
aud[18694]=16'hd8b5;
aud[18695]=16'hd8c6;
aud[18696]=16'hd8d7;
aud[18697]=16'hd8e8;
aud[18698]=16'hd8f9;
aud[18699]=16'hd90a;
aud[18700]=16'hd91b;
aud[18701]=16'hd92c;
aud[18702]=16'hd93d;
aud[18703]=16'hd94e;
aud[18704]=16'hd95f;
aud[18705]=16'hd970;
aud[18706]=16'hd982;
aud[18707]=16'hd993;
aud[18708]=16'hd9a4;
aud[18709]=16'hd9b5;
aud[18710]=16'hd9c6;
aud[18711]=16'hd9d7;
aud[18712]=16'hd9e9;
aud[18713]=16'hd9fa;
aud[18714]=16'hda0b;
aud[18715]=16'hda1c;
aud[18716]=16'hda2e;
aud[18717]=16'hda3f;
aud[18718]=16'hda50;
aud[18719]=16'hda62;
aud[18720]=16'hda73;
aud[18721]=16'hda84;
aud[18722]=16'hda96;
aud[18723]=16'hdaa7;
aud[18724]=16'hdab9;
aud[18725]=16'hdaca;
aud[18726]=16'hdadc;
aud[18727]=16'hdaed;
aud[18728]=16'hdaff;
aud[18729]=16'hdb10;
aud[18730]=16'hdb22;
aud[18731]=16'hdb33;
aud[18732]=16'hdb45;
aud[18733]=16'hdb56;
aud[18734]=16'hdb68;
aud[18735]=16'hdb79;
aud[18736]=16'hdb8b;
aud[18737]=16'hdb9d;
aud[18738]=16'hdbae;
aud[18739]=16'hdbc0;
aud[18740]=16'hdbd2;
aud[18741]=16'hdbe3;
aud[18742]=16'hdbf5;
aud[18743]=16'hdc07;
aud[18744]=16'hdc19;
aud[18745]=16'hdc2a;
aud[18746]=16'hdc3c;
aud[18747]=16'hdc4e;
aud[18748]=16'hdc60;
aud[18749]=16'hdc72;
aud[18750]=16'hdc83;
aud[18751]=16'hdc95;
aud[18752]=16'hdca7;
aud[18753]=16'hdcb9;
aud[18754]=16'hdccb;
aud[18755]=16'hdcdd;
aud[18756]=16'hdcef;
aud[18757]=16'hdd01;
aud[18758]=16'hdd13;
aud[18759]=16'hdd25;
aud[18760]=16'hdd37;
aud[18761]=16'hdd49;
aud[18762]=16'hdd5b;
aud[18763]=16'hdd6d;
aud[18764]=16'hdd7f;
aud[18765]=16'hdd91;
aud[18766]=16'hdda3;
aud[18767]=16'hddb5;
aud[18768]=16'hddc7;
aud[18769]=16'hddd9;
aud[18770]=16'hddeb;
aud[18771]=16'hddfe;
aud[18772]=16'hde10;
aud[18773]=16'hde22;
aud[18774]=16'hde34;
aud[18775]=16'hde46;
aud[18776]=16'hde59;
aud[18777]=16'hde6b;
aud[18778]=16'hde7d;
aud[18779]=16'hde8f;
aud[18780]=16'hdea2;
aud[18781]=16'hdeb4;
aud[18782]=16'hdec6;
aud[18783]=16'hded9;
aud[18784]=16'hdeeb;
aud[18785]=16'hdefd;
aud[18786]=16'hdf10;
aud[18787]=16'hdf22;
aud[18788]=16'hdf35;
aud[18789]=16'hdf47;
aud[18790]=16'hdf59;
aud[18791]=16'hdf6c;
aud[18792]=16'hdf7e;
aud[18793]=16'hdf91;
aud[18794]=16'hdfa3;
aud[18795]=16'hdfb6;
aud[18796]=16'hdfc8;
aud[18797]=16'hdfdb;
aud[18798]=16'hdfed;
aud[18799]=16'he000;
aud[18800]=16'he013;
aud[18801]=16'he025;
aud[18802]=16'he038;
aud[18803]=16'he04a;
aud[18804]=16'he05d;
aud[18805]=16'he070;
aud[18806]=16'he082;
aud[18807]=16'he095;
aud[18808]=16'he0a8;
aud[18809]=16'he0ba;
aud[18810]=16'he0cd;
aud[18811]=16'he0e0;
aud[18812]=16'he0f3;
aud[18813]=16'he105;
aud[18814]=16'he118;
aud[18815]=16'he12b;
aud[18816]=16'he13e;
aud[18817]=16'he151;
aud[18818]=16'he163;
aud[18819]=16'he176;
aud[18820]=16'he189;
aud[18821]=16'he19c;
aud[18822]=16'he1af;
aud[18823]=16'he1c2;
aud[18824]=16'he1d5;
aud[18825]=16'he1e8;
aud[18826]=16'he1fa;
aud[18827]=16'he20d;
aud[18828]=16'he220;
aud[18829]=16'he233;
aud[18830]=16'he246;
aud[18831]=16'he259;
aud[18832]=16'he26c;
aud[18833]=16'he27f;
aud[18834]=16'he292;
aud[18835]=16'he2a5;
aud[18836]=16'he2b9;
aud[18837]=16'he2cc;
aud[18838]=16'he2df;
aud[18839]=16'he2f2;
aud[18840]=16'he305;
aud[18841]=16'he318;
aud[18842]=16'he32b;
aud[18843]=16'he33e;
aud[18844]=16'he352;
aud[18845]=16'he365;
aud[18846]=16'he378;
aud[18847]=16'he38b;
aud[18848]=16'he39e;
aud[18849]=16'he3b2;
aud[18850]=16'he3c5;
aud[18851]=16'he3d8;
aud[18852]=16'he3eb;
aud[18853]=16'he3ff;
aud[18854]=16'he412;
aud[18855]=16'he425;
aud[18856]=16'he438;
aud[18857]=16'he44c;
aud[18858]=16'he45f;
aud[18859]=16'he473;
aud[18860]=16'he486;
aud[18861]=16'he499;
aud[18862]=16'he4ad;
aud[18863]=16'he4c0;
aud[18864]=16'he4d3;
aud[18865]=16'he4e7;
aud[18866]=16'he4fa;
aud[18867]=16'he50e;
aud[18868]=16'he521;
aud[18869]=16'he535;
aud[18870]=16'he548;
aud[18871]=16'he55c;
aud[18872]=16'he56f;
aud[18873]=16'he583;
aud[18874]=16'he596;
aud[18875]=16'he5aa;
aud[18876]=16'he5bd;
aud[18877]=16'he5d1;
aud[18878]=16'he5e4;
aud[18879]=16'he5f8;
aud[18880]=16'he60c;
aud[18881]=16'he61f;
aud[18882]=16'he633;
aud[18883]=16'he646;
aud[18884]=16'he65a;
aud[18885]=16'he66e;
aud[18886]=16'he681;
aud[18887]=16'he695;
aud[18888]=16'he6a9;
aud[18889]=16'he6bd;
aud[18890]=16'he6d0;
aud[18891]=16'he6e4;
aud[18892]=16'he6f8;
aud[18893]=16'he70b;
aud[18894]=16'he71f;
aud[18895]=16'he733;
aud[18896]=16'he747;
aud[18897]=16'he75b;
aud[18898]=16'he76e;
aud[18899]=16'he782;
aud[18900]=16'he796;
aud[18901]=16'he7aa;
aud[18902]=16'he7be;
aud[18903]=16'he7d1;
aud[18904]=16'he7e5;
aud[18905]=16'he7f9;
aud[18906]=16'he80d;
aud[18907]=16'he821;
aud[18908]=16'he835;
aud[18909]=16'he849;
aud[18910]=16'he85d;
aud[18911]=16'he871;
aud[18912]=16'he885;
aud[18913]=16'he899;
aud[18914]=16'he8ad;
aud[18915]=16'he8c0;
aud[18916]=16'he8d4;
aud[18917]=16'he8e8;
aud[18918]=16'he8fc;
aud[18919]=16'he910;
aud[18920]=16'he925;
aud[18921]=16'he939;
aud[18922]=16'he94d;
aud[18923]=16'he961;
aud[18924]=16'he975;
aud[18925]=16'he989;
aud[18926]=16'he99d;
aud[18927]=16'he9b1;
aud[18928]=16'he9c5;
aud[18929]=16'he9d9;
aud[18930]=16'he9ed;
aud[18931]=16'hea01;
aud[18932]=16'hea16;
aud[18933]=16'hea2a;
aud[18934]=16'hea3e;
aud[18935]=16'hea52;
aud[18936]=16'hea66;
aud[18937]=16'hea7a;
aud[18938]=16'hea8f;
aud[18939]=16'heaa3;
aud[18940]=16'heab7;
aud[18941]=16'heacb;
aud[18942]=16'heae0;
aud[18943]=16'heaf4;
aud[18944]=16'heb08;
aud[18945]=16'heb1c;
aud[18946]=16'heb31;
aud[18947]=16'heb45;
aud[18948]=16'heb59;
aud[18949]=16'heb6e;
aud[18950]=16'heb82;
aud[18951]=16'heb96;
aud[18952]=16'hebab;
aud[18953]=16'hebbf;
aud[18954]=16'hebd3;
aud[18955]=16'hebe8;
aud[18956]=16'hebfc;
aud[18957]=16'hec10;
aud[18958]=16'hec25;
aud[18959]=16'hec39;
aud[18960]=16'hec4d;
aud[18961]=16'hec62;
aud[18962]=16'hec76;
aud[18963]=16'hec8b;
aud[18964]=16'hec9f;
aud[18965]=16'hecb4;
aud[18966]=16'hecc8;
aud[18967]=16'hecdd;
aud[18968]=16'hecf1;
aud[18969]=16'hed05;
aud[18970]=16'hed1a;
aud[18971]=16'hed2e;
aud[18972]=16'hed43;
aud[18973]=16'hed57;
aud[18974]=16'hed6c;
aud[18975]=16'hed81;
aud[18976]=16'hed95;
aud[18977]=16'hedaa;
aud[18978]=16'hedbe;
aud[18979]=16'hedd3;
aud[18980]=16'hede7;
aud[18981]=16'hedfc;
aud[18982]=16'hee10;
aud[18983]=16'hee25;
aud[18984]=16'hee3a;
aud[18985]=16'hee4e;
aud[18986]=16'hee63;
aud[18987]=16'hee77;
aud[18988]=16'hee8c;
aud[18989]=16'heea1;
aud[18990]=16'heeb5;
aud[18991]=16'heeca;
aud[18992]=16'heedf;
aud[18993]=16'heef3;
aud[18994]=16'hef08;
aud[18995]=16'hef1d;
aud[18996]=16'hef31;
aud[18997]=16'hef46;
aud[18998]=16'hef5b;
aud[18999]=16'hef70;
aud[19000]=16'hef84;
aud[19001]=16'hef99;
aud[19002]=16'hefae;
aud[19003]=16'hefc2;
aud[19004]=16'hefd7;
aud[19005]=16'hefec;
aud[19006]=16'hf001;
aud[19007]=16'hf015;
aud[19008]=16'hf02a;
aud[19009]=16'hf03f;
aud[19010]=16'hf054;
aud[19011]=16'hf069;
aud[19012]=16'hf07d;
aud[19013]=16'hf092;
aud[19014]=16'hf0a7;
aud[19015]=16'hf0bc;
aud[19016]=16'hf0d1;
aud[19017]=16'hf0e6;
aud[19018]=16'hf0fa;
aud[19019]=16'hf10f;
aud[19020]=16'hf124;
aud[19021]=16'hf139;
aud[19022]=16'hf14e;
aud[19023]=16'hf163;
aud[19024]=16'hf178;
aud[19025]=16'hf18c;
aud[19026]=16'hf1a1;
aud[19027]=16'hf1b6;
aud[19028]=16'hf1cb;
aud[19029]=16'hf1e0;
aud[19030]=16'hf1f5;
aud[19031]=16'hf20a;
aud[19032]=16'hf21f;
aud[19033]=16'hf234;
aud[19034]=16'hf249;
aud[19035]=16'hf25e;
aud[19036]=16'hf273;
aud[19037]=16'hf288;
aud[19038]=16'hf29d;
aud[19039]=16'hf2b2;
aud[19040]=16'hf2c7;
aud[19041]=16'hf2dc;
aud[19042]=16'hf2f1;
aud[19043]=16'hf306;
aud[19044]=16'hf31b;
aud[19045]=16'hf330;
aud[19046]=16'hf345;
aud[19047]=16'hf35a;
aud[19048]=16'hf36f;
aud[19049]=16'hf384;
aud[19050]=16'hf399;
aud[19051]=16'hf3ae;
aud[19052]=16'hf3c3;
aud[19053]=16'hf3d8;
aud[19054]=16'hf3ed;
aud[19055]=16'hf402;
aud[19056]=16'hf417;
aud[19057]=16'hf42c;
aud[19058]=16'hf441;
aud[19059]=16'hf456;
aud[19060]=16'hf46b;
aud[19061]=16'hf480;
aud[19062]=16'hf496;
aud[19063]=16'hf4ab;
aud[19064]=16'hf4c0;
aud[19065]=16'hf4d5;
aud[19066]=16'hf4ea;
aud[19067]=16'hf4ff;
aud[19068]=16'hf514;
aud[19069]=16'hf529;
aud[19070]=16'hf53f;
aud[19071]=16'hf554;
aud[19072]=16'hf569;
aud[19073]=16'hf57e;
aud[19074]=16'hf593;
aud[19075]=16'hf5a8;
aud[19076]=16'hf5bd;
aud[19077]=16'hf5d3;
aud[19078]=16'hf5e8;
aud[19079]=16'hf5fd;
aud[19080]=16'hf612;
aud[19081]=16'hf627;
aud[19082]=16'hf63d;
aud[19083]=16'hf652;
aud[19084]=16'hf667;
aud[19085]=16'hf67c;
aud[19086]=16'hf691;
aud[19087]=16'hf6a7;
aud[19088]=16'hf6bc;
aud[19089]=16'hf6d1;
aud[19090]=16'hf6e6;
aud[19091]=16'hf6fb;
aud[19092]=16'hf711;
aud[19093]=16'hf726;
aud[19094]=16'hf73b;
aud[19095]=16'hf750;
aud[19096]=16'hf766;
aud[19097]=16'hf77b;
aud[19098]=16'hf790;
aud[19099]=16'hf7a5;
aud[19100]=16'hf7bb;
aud[19101]=16'hf7d0;
aud[19102]=16'hf7e5;
aud[19103]=16'hf7fb;
aud[19104]=16'hf810;
aud[19105]=16'hf825;
aud[19106]=16'hf83a;
aud[19107]=16'hf850;
aud[19108]=16'hf865;
aud[19109]=16'hf87a;
aud[19110]=16'hf890;
aud[19111]=16'hf8a5;
aud[19112]=16'hf8ba;
aud[19113]=16'hf8cf;
aud[19114]=16'hf8e5;
aud[19115]=16'hf8fa;
aud[19116]=16'hf90f;
aud[19117]=16'hf925;
aud[19118]=16'hf93a;
aud[19119]=16'hf94f;
aud[19120]=16'hf965;
aud[19121]=16'hf97a;
aud[19122]=16'hf98f;
aud[19123]=16'hf9a5;
aud[19124]=16'hf9ba;
aud[19125]=16'hf9cf;
aud[19126]=16'hf9e5;
aud[19127]=16'hf9fa;
aud[19128]=16'hfa0f;
aud[19129]=16'hfa25;
aud[19130]=16'hfa3a;
aud[19131]=16'hfa50;
aud[19132]=16'hfa65;
aud[19133]=16'hfa7a;
aud[19134]=16'hfa90;
aud[19135]=16'hfaa5;
aud[19136]=16'hfaba;
aud[19137]=16'hfad0;
aud[19138]=16'hfae5;
aud[19139]=16'hfafb;
aud[19140]=16'hfb10;
aud[19141]=16'hfb25;
aud[19142]=16'hfb3b;
aud[19143]=16'hfb50;
aud[19144]=16'hfb65;
aud[19145]=16'hfb7b;
aud[19146]=16'hfb90;
aud[19147]=16'hfba6;
aud[19148]=16'hfbbb;
aud[19149]=16'hfbd0;
aud[19150]=16'hfbe6;
aud[19151]=16'hfbfb;
aud[19152]=16'hfc11;
aud[19153]=16'hfc26;
aud[19154]=16'hfc3b;
aud[19155]=16'hfc51;
aud[19156]=16'hfc66;
aud[19157]=16'hfc7c;
aud[19158]=16'hfc91;
aud[19159]=16'hfca7;
aud[19160]=16'hfcbc;
aud[19161]=16'hfcd1;
aud[19162]=16'hfce7;
aud[19163]=16'hfcfc;
aud[19164]=16'hfd12;
aud[19165]=16'hfd27;
aud[19166]=16'hfd3c;
aud[19167]=16'hfd52;
aud[19168]=16'hfd67;
aud[19169]=16'hfd7d;
aud[19170]=16'hfd92;
aud[19171]=16'hfda8;
aud[19172]=16'hfdbd;
aud[19173]=16'hfdd2;
aud[19174]=16'hfde8;
aud[19175]=16'hfdfd;
aud[19176]=16'hfe13;
aud[19177]=16'hfe28;
aud[19178]=16'hfe3e;
aud[19179]=16'hfe53;
aud[19180]=16'hfe69;
aud[19181]=16'hfe7e;
aud[19182]=16'hfe93;
aud[19183]=16'hfea9;
aud[19184]=16'hfebe;
aud[19185]=16'hfed4;
aud[19186]=16'hfee9;
aud[19187]=16'hfeff;
aud[19188]=16'hff14;
aud[19189]=16'hff2a;
aud[19190]=16'hff3f;
aud[19191]=16'hff54;
aud[19192]=16'hff6a;
aud[19193]=16'hff7f;
aud[19194]=16'hff95;
aud[19195]=16'hffaa;
aud[19196]=16'hffc0;
aud[19197]=16'hffd5;
aud[19198]=16'hffeb;
aud[19199]=16'h0;
aud[19200]=16'h15;
aud[19201]=16'h2b;
aud[19202]=16'h40;
aud[19203]=16'h56;
aud[19204]=16'h6b;
aud[19205]=16'h81;
aud[19206]=16'h96;
aud[19207]=16'hac;
aud[19208]=16'hc1;
aud[19209]=16'hd6;
aud[19210]=16'hec;
aud[19211]=16'h101;
aud[19212]=16'h117;
aud[19213]=16'h12c;
aud[19214]=16'h142;
aud[19215]=16'h157;
aud[19216]=16'h16d;
aud[19217]=16'h182;
aud[19218]=16'h197;
aud[19219]=16'h1ad;
aud[19220]=16'h1c2;
aud[19221]=16'h1d8;
aud[19222]=16'h1ed;
aud[19223]=16'h203;
aud[19224]=16'h218;
aud[19225]=16'h22e;
aud[19226]=16'h243;
aud[19227]=16'h258;
aud[19228]=16'h26e;
aud[19229]=16'h283;
aud[19230]=16'h299;
aud[19231]=16'h2ae;
aud[19232]=16'h2c4;
aud[19233]=16'h2d9;
aud[19234]=16'h2ee;
aud[19235]=16'h304;
aud[19236]=16'h319;
aud[19237]=16'h32f;
aud[19238]=16'h344;
aud[19239]=16'h359;
aud[19240]=16'h36f;
aud[19241]=16'h384;
aud[19242]=16'h39a;
aud[19243]=16'h3af;
aud[19244]=16'h3c5;
aud[19245]=16'h3da;
aud[19246]=16'h3ef;
aud[19247]=16'h405;
aud[19248]=16'h41a;
aud[19249]=16'h430;
aud[19250]=16'h445;
aud[19251]=16'h45a;
aud[19252]=16'h470;
aud[19253]=16'h485;
aud[19254]=16'h49b;
aud[19255]=16'h4b0;
aud[19256]=16'h4c5;
aud[19257]=16'h4db;
aud[19258]=16'h4f0;
aud[19259]=16'h505;
aud[19260]=16'h51b;
aud[19261]=16'h530;
aud[19262]=16'h546;
aud[19263]=16'h55b;
aud[19264]=16'h570;
aud[19265]=16'h586;
aud[19266]=16'h59b;
aud[19267]=16'h5b0;
aud[19268]=16'h5c6;
aud[19269]=16'h5db;
aud[19270]=16'h5f1;
aud[19271]=16'h606;
aud[19272]=16'h61b;
aud[19273]=16'h631;
aud[19274]=16'h646;
aud[19275]=16'h65b;
aud[19276]=16'h671;
aud[19277]=16'h686;
aud[19278]=16'h69b;
aud[19279]=16'h6b1;
aud[19280]=16'h6c6;
aud[19281]=16'h6db;
aud[19282]=16'h6f1;
aud[19283]=16'h706;
aud[19284]=16'h71b;
aud[19285]=16'h731;
aud[19286]=16'h746;
aud[19287]=16'h75b;
aud[19288]=16'h770;
aud[19289]=16'h786;
aud[19290]=16'h79b;
aud[19291]=16'h7b0;
aud[19292]=16'h7c6;
aud[19293]=16'h7db;
aud[19294]=16'h7f0;
aud[19295]=16'h805;
aud[19296]=16'h81b;
aud[19297]=16'h830;
aud[19298]=16'h845;
aud[19299]=16'h85b;
aud[19300]=16'h870;
aud[19301]=16'h885;
aud[19302]=16'h89a;
aud[19303]=16'h8b0;
aud[19304]=16'h8c5;
aud[19305]=16'h8da;
aud[19306]=16'h8ef;
aud[19307]=16'h905;
aud[19308]=16'h91a;
aud[19309]=16'h92f;
aud[19310]=16'h944;
aud[19311]=16'h959;
aud[19312]=16'h96f;
aud[19313]=16'h984;
aud[19314]=16'h999;
aud[19315]=16'h9ae;
aud[19316]=16'h9c3;
aud[19317]=16'h9d9;
aud[19318]=16'h9ee;
aud[19319]=16'ha03;
aud[19320]=16'ha18;
aud[19321]=16'ha2d;
aud[19322]=16'ha43;
aud[19323]=16'ha58;
aud[19324]=16'ha6d;
aud[19325]=16'ha82;
aud[19326]=16'ha97;
aud[19327]=16'haac;
aud[19328]=16'hac1;
aud[19329]=16'had7;
aud[19330]=16'haec;
aud[19331]=16'hb01;
aud[19332]=16'hb16;
aud[19333]=16'hb2b;
aud[19334]=16'hb40;
aud[19335]=16'hb55;
aud[19336]=16'hb6a;
aud[19337]=16'hb80;
aud[19338]=16'hb95;
aud[19339]=16'hbaa;
aud[19340]=16'hbbf;
aud[19341]=16'hbd4;
aud[19342]=16'hbe9;
aud[19343]=16'hbfe;
aud[19344]=16'hc13;
aud[19345]=16'hc28;
aud[19346]=16'hc3d;
aud[19347]=16'hc52;
aud[19348]=16'hc67;
aud[19349]=16'hc7c;
aud[19350]=16'hc91;
aud[19351]=16'hca6;
aud[19352]=16'hcbb;
aud[19353]=16'hcd0;
aud[19354]=16'hce5;
aud[19355]=16'hcfa;
aud[19356]=16'hd0f;
aud[19357]=16'hd24;
aud[19358]=16'hd39;
aud[19359]=16'hd4e;
aud[19360]=16'hd63;
aud[19361]=16'hd78;
aud[19362]=16'hd8d;
aud[19363]=16'hda2;
aud[19364]=16'hdb7;
aud[19365]=16'hdcc;
aud[19366]=16'hde1;
aud[19367]=16'hdf6;
aud[19368]=16'he0b;
aud[19369]=16'he20;
aud[19370]=16'he35;
aud[19371]=16'he4a;
aud[19372]=16'he5f;
aud[19373]=16'he74;
aud[19374]=16'he88;
aud[19375]=16'he9d;
aud[19376]=16'heb2;
aud[19377]=16'hec7;
aud[19378]=16'hedc;
aud[19379]=16'hef1;
aud[19380]=16'hf06;
aud[19381]=16'hf1a;
aud[19382]=16'hf2f;
aud[19383]=16'hf44;
aud[19384]=16'hf59;
aud[19385]=16'hf6e;
aud[19386]=16'hf83;
aud[19387]=16'hf97;
aud[19388]=16'hfac;
aud[19389]=16'hfc1;
aud[19390]=16'hfd6;
aud[19391]=16'hfeb;
aud[19392]=16'hfff;
aud[19393]=16'h1014;
aud[19394]=16'h1029;
aud[19395]=16'h103e;
aud[19396]=16'h1052;
aud[19397]=16'h1067;
aud[19398]=16'h107c;
aud[19399]=16'h1090;
aud[19400]=16'h10a5;
aud[19401]=16'h10ba;
aud[19402]=16'h10cf;
aud[19403]=16'h10e3;
aud[19404]=16'h10f8;
aud[19405]=16'h110d;
aud[19406]=16'h1121;
aud[19407]=16'h1136;
aud[19408]=16'h114b;
aud[19409]=16'h115f;
aud[19410]=16'h1174;
aud[19411]=16'h1189;
aud[19412]=16'h119d;
aud[19413]=16'h11b2;
aud[19414]=16'h11c6;
aud[19415]=16'h11db;
aud[19416]=16'h11f0;
aud[19417]=16'h1204;
aud[19418]=16'h1219;
aud[19419]=16'h122d;
aud[19420]=16'h1242;
aud[19421]=16'h1256;
aud[19422]=16'h126b;
aud[19423]=16'h127f;
aud[19424]=16'h1294;
aud[19425]=16'h12a9;
aud[19426]=16'h12bd;
aud[19427]=16'h12d2;
aud[19428]=16'h12e6;
aud[19429]=16'h12fb;
aud[19430]=16'h130f;
aud[19431]=16'h1323;
aud[19432]=16'h1338;
aud[19433]=16'h134c;
aud[19434]=16'h1361;
aud[19435]=16'h1375;
aud[19436]=16'h138a;
aud[19437]=16'h139e;
aud[19438]=16'h13b3;
aud[19439]=16'h13c7;
aud[19440]=16'h13db;
aud[19441]=16'h13f0;
aud[19442]=16'h1404;
aud[19443]=16'h1418;
aud[19444]=16'h142d;
aud[19445]=16'h1441;
aud[19446]=16'h1455;
aud[19447]=16'h146a;
aud[19448]=16'h147e;
aud[19449]=16'h1492;
aud[19450]=16'h14a7;
aud[19451]=16'h14bb;
aud[19452]=16'h14cf;
aud[19453]=16'h14e4;
aud[19454]=16'h14f8;
aud[19455]=16'h150c;
aud[19456]=16'h1520;
aud[19457]=16'h1535;
aud[19458]=16'h1549;
aud[19459]=16'h155d;
aud[19460]=16'h1571;
aud[19461]=16'h1586;
aud[19462]=16'h159a;
aud[19463]=16'h15ae;
aud[19464]=16'h15c2;
aud[19465]=16'h15d6;
aud[19466]=16'h15ea;
aud[19467]=16'h15ff;
aud[19468]=16'h1613;
aud[19469]=16'h1627;
aud[19470]=16'h163b;
aud[19471]=16'h164f;
aud[19472]=16'h1663;
aud[19473]=16'h1677;
aud[19474]=16'h168b;
aud[19475]=16'h169f;
aud[19476]=16'h16b3;
aud[19477]=16'h16c7;
aud[19478]=16'h16db;
aud[19479]=16'h16f0;
aud[19480]=16'h1704;
aud[19481]=16'h1718;
aud[19482]=16'h172c;
aud[19483]=16'h1740;
aud[19484]=16'h1753;
aud[19485]=16'h1767;
aud[19486]=16'h177b;
aud[19487]=16'h178f;
aud[19488]=16'h17a3;
aud[19489]=16'h17b7;
aud[19490]=16'h17cb;
aud[19491]=16'h17df;
aud[19492]=16'h17f3;
aud[19493]=16'h1807;
aud[19494]=16'h181b;
aud[19495]=16'h182f;
aud[19496]=16'h1842;
aud[19497]=16'h1856;
aud[19498]=16'h186a;
aud[19499]=16'h187e;
aud[19500]=16'h1892;
aud[19501]=16'h18a5;
aud[19502]=16'h18b9;
aud[19503]=16'h18cd;
aud[19504]=16'h18e1;
aud[19505]=16'h18f5;
aud[19506]=16'h1908;
aud[19507]=16'h191c;
aud[19508]=16'h1930;
aud[19509]=16'h1943;
aud[19510]=16'h1957;
aud[19511]=16'h196b;
aud[19512]=16'h197f;
aud[19513]=16'h1992;
aud[19514]=16'h19a6;
aud[19515]=16'h19ba;
aud[19516]=16'h19cd;
aud[19517]=16'h19e1;
aud[19518]=16'h19f4;
aud[19519]=16'h1a08;
aud[19520]=16'h1a1c;
aud[19521]=16'h1a2f;
aud[19522]=16'h1a43;
aud[19523]=16'h1a56;
aud[19524]=16'h1a6a;
aud[19525]=16'h1a7d;
aud[19526]=16'h1a91;
aud[19527]=16'h1aa4;
aud[19528]=16'h1ab8;
aud[19529]=16'h1acb;
aud[19530]=16'h1adf;
aud[19531]=16'h1af2;
aud[19532]=16'h1b06;
aud[19533]=16'h1b19;
aud[19534]=16'h1b2d;
aud[19535]=16'h1b40;
aud[19536]=16'h1b53;
aud[19537]=16'h1b67;
aud[19538]=16'h1b7a;
aud[19539]=16'h1b8d;
aud[19540]=16'h1ba1;
aud[19541]=16'h1bb4;
aud[19542]=16'h1bc8;
aud[19543]=16'h1bdb;
aud[19544]=16'h1bee;
aud[19545]=16'h1c01;
aud[19546]=16'h1c15;
aud[19547]=16'h1c28;
aud[19548]=16'h1c3b;
aud[19549]=16'h1c4e;
aud[19550]=16'h1c62;
aud[19551]=16'h1c75;
aud[19552]=16'h1c88;
aud[19553]=16'h1c9b;
aud[19554]=16'h1cae;
aud[19555]=16'h1cc2;
aud[19556]=16'h1cd5;
aud[19557]=16'h1ce8;
aud[19558]=16'h1cfb;
aud[19559]=16'h1d0e;
aud[19560]=16'h1d21;
aud[19561]=16'h1d34;
aud[19562]=16'h1d47;
aud[19563]=16'h1d5b;
aud[19564]=16'h1d6e;
aud[19565]=16'h1d81;
aud[19566]=16'h1d94;
aud[19567]=16'h1da7;
aud[19568]=16'h1dba;
aud[19569]=16'h1dcd;
aud[19570]=16'h1de0;
aud[19571]=16'h1df3;
aud[19572]=16'h1e06;
aud[19573]=16'h1e18;
aud[19574]=16'h1e2b;
aud[19575]=16'h1e3e;
aud[19576]=16'h1e51;
aud[19577]=16'h1e64;
aud[19578]=16'h1e77;
aud[19579]=16'h1e8a;
aud[19580]=16'h1e9d;
aud[19581]=16'h1eaf;
aud[19582]=16'h1ec2;
aud[19583]=16'h1ed5;
aud[19584]=16'h1ee8;
aud[19585]=16'h1efb;
aud[19586]=16'h1f0d;
aud[19587]=16'h1f20;
aud[19588]=16'h1f33;
aud[19589]=16'h1f46;
aud[19590]=16'h1f58;
aud[19591]=16'h1f6b;
aud[19592]=16'h1f7e;
aud[19593]=16'h1f90;
aud[19594]=16'h1fa3;
aud[19595]=16'h1fb6;
aud[19596]=16'h1fc8;
aud[19597]=16'h1fdb;
aud[19598]=16'h1fed;
aud[19599]=16'h2000;
aud[19600]=16'h2013;
aud[19601]=16'h2025;
aud[19602]=16'h2038;
aud[19603]=16'h204a;
aud[19604]=16'h205d;
aud[19605]=16'h206f;
aud[19606]=16'h2082;
aud[19607]=16'h2094;
aud[19608]=16'h20a7;
aud[19609]=16'h20b9;
aud[19610]=16'h20cb;
aud[19611]=16'h20de;
aud[19612]=16'h20f0;
aud[19613]=16'h2103;
aud[19614]=16'h2115;
aud[19615]=16'h2127;
aud[19616]=16'h213a;
aud[19617]=16'h214c;
aud[19618]=16'h215e;
aud[19619]=16'h2171;
aud[19620]=16'h2183;
aud[19621]=16'h2195;
aud[19622]=16'h21a7;
aud[19623]=16'h21ba;
aud[19624]=16'h21cc;
aud[19625]=16'h21de;
aud[19626]=16'h21f0;
aud[19627]=16'h2202;
aud[19628]=16'h2215;
aud[19629]=16'h2227;
aud[19630]=16'h2239;
aud[19631]=16'h224b;
aud[19632]=16'h225d;
aud[19633]=16'h226f;
aud[19634]=16'h2281;
aud[19635]=16'h2293;
aud[19636]=16'h22a5;
aud[19637]=16'h22b7;
aud[19638]=16'h22c9;
aud[19639]=16'h22db;
aud[19640]=16'h22ed;
aud[19641]=16'h22ff;
aud[19642]=16'h2311;
aud[19643]=16'h2323;
aud[19644]=16'h2335;
aud[19645]=16'h2347;
aud[19646]=16'h2359;
aud[19647]=16'h236b;
aud[19648]=16'h237d;
aud[19649]=16'h238e;
aud[19650]=16'h23a0;
aud[19651]=16'h23b2;
aud[19652]=16'h23c4;
aud[19653]=16'h23d6;
aud[19654]=16'h23e7;
aud[19655]=16'h23f9;
aud[19656]=16'h240b;
aud[19657]=16'h241d;
aud[19658]=16'h242e;
aud[19659]=16'h2440;
aud[19660]=16'h2452;
aud[19661]=16'h2463;
aud[19662]=16'h2475;
aud[19663]=16'h2487;
aud[19664]=16'h2498;
aud[19665]=16'h24aa;
aud[19666]=16'h24bb;
aud[19667]=16'h24cd;
aud[19668]=16'h24de;
aud[19669]=16'h24f0;
aud[19670]=16'h2501;
aud[19671]=16'h2513;
aud[19672]=16'h2524;
aud[19673]=16'h2536;
aud[19674]=16'h2547;
aud[19675]=16'h2559;
aud[19676]=16'h256a;
aud[19677]=16'h257c;
aud[19678]=16'h258d;
aud[19679]=16'h259e;
aud[19680]=16'h25b0;
aud[19681]=16'h25c1;
aud[19682]=16'h25d2;
aud[19683]=16'h25e4;
aud[19684]=16'h25f5;
aud[19685]=16'h2606;
aud[19686]=16'h2617;
aud[19687]=16'h2629;
aud[19688]=16'h263a;
aud[19689]=16'h264b;
aud[19690]=16'h265c;
aud[19691]=16'h266d;
aud[19692]=16'h267e;
aud[19693]=16'h2690;
aud[19694]=16'h26a1;
aud[19695]=16'h26b2;
aud[19696]=16'h26c3;
aud[19697]=16'h26d4;
aud[19698]=16'h26e5;
aud[19699]=16'h26f6;
aud[19700]=16'h2707;
aud[19701]=16'h2718;
aud[19702]=16'h2729;
aud[19703]=16'h273a;
aud[19704]=16'h274b;
aud[19705]=16'h275c;
aud[19706]=16'h276d;
aud[19707]=16'h277e;
aud[19708]=16'h278e;
aud[19709]=16'h279f;
aud[19710]=16'h27b0;
aud[19711]=16'h27c1;
aud[19712]=16'h27d2;
aud[19713]=16'h27e2;
aud[19714]=16'h27f3;
aud[19715]=16'h2804;
aud[19716]=16'h2815;
aud[19717]=16'h2825;
aud[19718]=16'h2836;
aud[19719]=16'h2847;
aud[19720]=16'h2857;
aud[19721]=16'h2868;
aud[19722]=16'h2879;
aud[19723]=16'h2889;
aud[19724]=16'h289a;
aud[19725]=16'h28aa;
aud[19726]=16'h28bb;
aud[19727]=16'h28cc;
aud[19728]=16'h28dc;
aud[19729]=16'h28ed;
aud[19730]=16'h28fd;
aud[19731]=16'h290e;
aud[19732]=16'h291e;
aud[19733]=16'h292e;
aud[19734]=16'h293f;
aud[19735]=16'h294f;
aud[19736]=16'h2960;
aud[19737]=16'h2970;
aud[19738]=16'h2980;
aud[19739]=16'h2991;
aud[19740]=16'h29a1;
aud[19741]=16'h29b1;
aud[19742]=16'h29c1;
aud[19743]=16'h29d2;
aud[19744]=16'h29e2;
aud[19745]=16'h29f2;
aud[19746]=16'h2a02;
aud[19747]=16'h2a12;
aud[19748]=16'h2a23;
aud[19749]=16'h2a33;
aud[19750]=16'h2a43;
aud[19751]=16'h2a53;
aud[19752]=16'h2a63;
aud[19753]=16'h2a73;
aud[19754]=16'h2a83;
aud[19755]=16'h2a93;
aud[19756]=16'h2aa3;
aud[19757]=16'h2ab3;
aud[19758]=16'h2ac3;
aud[19759]=16'h2ad3;
aud[19760]=16'h2ae3;
aud[19761]=16'h2af3;
aud[19762]=16'h2b03;
aud[19763]=16'h2b13;
aud[19764]=16'h2b22;
aud[19765]=16'h2b32;
aud[19766]=16'h2b42;
aud[19767]=16'h2b52;
aud[19768]=16'h2b62;
aud[19769]=16'h2b71;
aud[19770]=16'h2b81;
aud[19771]=16'h2b91;
aud[19772]=16'h2ba1;
aud[19773]=16'h2bb0;
aud[19774]=16'h2bc0;
aud[19775]=16'h2bd0;
aud[19776]=16'h2bdf;
aud[19777]=16'h2bef;
aud[19778]=16'h2bfe;
aud[19779]=16'h2c0e;
aud[19780]=16'h2c1e;
aud[19781]=16'h2c2d;
aud[19782]=16'h2c3d;
aud[19783]=16'h2c4c;
aud[19784]=16'h2c5c;
aud[19785]=16'h2c6b;
aud[19786]=16'h2c7a;
aud[19787]=16'h2c8a;
aud[19788]=16'h2c99;
aud[19789]=16'h2ca9;
aud[19790]=16'h2cb8;
aud[19791]=16'h2cc7;
aud[19792]=16'h2cd7;
aud[19793]=16'h2ce6;
aud[19794]=16'h2cf5;
aud[19795]=16'h2d04;
aud[19796]=16'h2d14;
aud[19797]=16'h2d23;
aud[19798]=16'h2d32;
aud[19799]=16'h2d41;
aud[19800]=16'h2d50;
aud[19801]=16'h2d60;
aud[19802]=16'h2d6f;
aud[19803]=16'h2d7e;
aud[19804]=16'h2d8d;
aud[19805]=16'h2d9c;
aud[19806]=16'h2dab;
aud[19807]=16'h2dba;
aud[19808]=16'h2dc9;
aud[19809]=16'h2dd8;
aud[19810]=16'h2de7;
aud[19811]=16'h2df6;
aud[19812]=16'h2e05;
aud[19813]=16'h2e14;
aud[19814]=16'h2e22;
aud[19815]=16'h2e31;
aud[19816]=16'h2e40;
aud[19817]=16'h2e4f;
aud[19818]=16'h2e5e;
aud[19819]=16'h2e6d;
aud[19820]=16'h2e7b;
aud[19821]=16'h2e8a;
aud[19822]=16'h2e99;
aud[19823]=16'h2ea7;
aud[19824]=16'h2eb6;
aud[19825]=16'h2ec5;
aud[19826]=16'h2ed3;
aud[19827]=16'h2ee2;
aud[19828]=16'h2ef1;
aud[19829]=16'h2eff;
aud[19830]=16'h2f0e;
aud[19831]=16'h2f1c;
aud[19832]=16'h2f2b;
aud[19833]=16'h2f39;
aud[19834]=16'h2f48;
aud[19835]=16'h2f56;
aud[19836]=16'h2f65;
aud[19837]=16'h2f73;
aud[19838]=16'h2f81;
aud[19839]=16'h2f90;
aud[19840]=16'h2f9e;
aud[19841]=16'h2fac;
aud[19842]=16'h2fbb;
aud[19843]=16'h2fc9;
aud[19844]=16'h2fd7;
aud[19845]=16'h2fe5;
aud[19846]=16'h2ff4;
aud[19847]=16'h3002;
aud[19848]=16'h3010;
aud[19849]=16'h301e;
aud[19850]=16'h302c;
aud[19851]=16'h303a;
aud[19852]=16'h3048;
aud[19853]=16'h3057;
aud[19854]=16'h3065;
aud[19855]=16'h3073;
aud[19856]=16'h3081;
aud[19857]=16'h308f;
aud[19858]=16'h309d;
aud[19859]=16'h30aa;
aud[19860]=16'h30b8;
aud[19861]=16'h30c6;
aud[19862]=16'h30d4;
aud[19863]=16'h30e2;
aud[19864]=16'h30f0;
aud[19865]=16'h30fe;
aud[19866]=16'h310b;
aud[19867]=16'h3119;
aud[19868]=16'h3127;
aud[19869]=16'h3135;
aud[19870]=16'h3142;
aud[19871]=16'h3150;
aud[19872]=16'h315e;
aud[19873]=16'h316b;
aud[19874]=16'h3179;
aud[19875]=16'h3187;
aud[19876]=16'h3194;
aud[19877]=16'h31a2;
aud[19878]=16'h31af;
aud[19879]=16'h31bd;
aud[19880]=16'h31ca;
aud[19881]=16'h31d8;
aud[19882]=16'h31e5;
aud[19883]=16'h31f3;
aud[19884]=16'h3200;
aud[19885]=16'h320d;
aud[19886]=16'h321b;
aud[19887]=16'h3228;
aud[19888]=16'h3235;
aud[19889]=16'h3243;
aud[19890]=16'h3250;
aud[19891]=16'h325d;
aud[19892]=16'h326a;
aud[19893]=16'h3278;
aud[19894]=16'h3285;
aud[19895]=16'h3292;
aud[19896]=16'h329f;
aud[19897]=16'h32ac;
aud[19898]=16'h32b9;
aud[19899]=16'h32c6;
aud[19900]=16'h32d3;
aud[19901]=16'h32e0;
aud[19902]=16'h32ed;
aud[19903]=16'h32fa;
aud[19904]=16'h3307;
aud[19905]=16'h3314;
aud[19906]=16'h3321;
aud[19907]=16'h332e;
aud[19908]=16'h333b;
aud[19909]=16'h3348;
aud[19910]=16'h3355;
aud[19911]=16'h3361;
aud[19912]=16'h336e;
aud[19913]=16'h337b;
aud[19914]=16'h3388;
aud[19915]=16'h3394;
aud[19916]=16'h33a1;
aud[19917]=16'h33ae;
aud[19918]=16'h33ba;
aud[19919]=16'h33c7;
aud[19920]=16'h33d4;
aud[19921]=16'h33e0;
aud[19922]=16'h33ed;
aud[19923]=16'h33f9;
aud[19924]=16'h3406;
aud[19925]=16'h3412;
aud[19926]=16'h341f;
aud[19927]=16'h342b;
aud[19928]=16'h3437;
aud[19929]=16'h3444;
aud[19930]=16'h3450;
aud[19931]=16'h345d;
aud[19932]=16'h3469;
aud[19933]=16'h3475;
aud[19934]=16'h3481;
aud[19935]=16'h348e;
aud[19936]=16'h349a;
aud[19937]=16'h34a6;
aud[19938]=16'h34b2;
aud[19939]=16'h34be;
aud[19940]=16'h34cb;
aud[19941]=16'h34d7;
aud[19942]=16'h34e3;
aud[19943]=16'h34ef;
aud[19944]=16'h34fb;
aud[19945]=16'h3507;
aud[19946]=16'h3513;
aud[19947]=16'h351f;
aud[19948]=16'h352b;
aud[19949]=16'h3537;
aud[19950]=16'h3543;
aud[19951]=16'h354f;
aud[19952]=16'h355a;
aud[19953]=16'h3566;
aud[19954]=16'h3572;
aud[19955]=16'h357e;
aud[19956]=16'h358a;
aud[19957]=16'h3595;
aud[19958]=16'h35a1;
aud[19959]=16'h35ad;
aud[19960]=16'h35b8;
aud[19961]=16'h35c4;
aud[19962]=16'h35d0;
aud[19963]=16'h35db;
aud[19964]=16'h35e7;
aud[19965]=16'h35f2;
aud[19966]=16'h35fe;
aud[19967]=16'h3609;
aud[19968]=16'h3615;
aud[19969]=16'h3620;
aud[19970]=16'h362c;
aud[19971]=16'h3637;
aud[19972]=16'h3643;
aud[19973]=16'h364e;
aud[19974]=16'h3659;
aud[19975]=16'h3665;
aud[19976]=16'h3670;
aud[19977]=16'h367b;
aud[19978]=16'h3686;
aud[19979]=16'h3692;
aud[19980]=16'h369d;
aud[19981]=16'h36a8;
aud[19982]=16'h36b3;
aud[19983]=16'h36be;
aud[19984]=16'h36c9;
aud[19985]=16'h36d4;
aud[19986]=16'h36e0;
aud[19987]=16'h36eb;
aud[19988]=16'h36f6;
aud[19989]=16'h3701;
aud[19990]=16'h370b;
aud[19991]=16'h3716;
aud[19992]=16'h3721;
aud[19993]=16'h372c;
aud[19994]=16'h3737;
aud[19995]=16'h3742;
aud[19996]=16'h374d;
aud[19997]=16'h3757;
aud[19998]=16'h3762;
aud[19999]=16'h376d;
aud[20000]=16'h3778;
aud[20001]=16'h3782;
aud[20002]=16'h378d;
aud[20003]=16'h3798;
aud[20004]=16'h37a2;
aud[20005]=16'h37ad;
aud[20006]=16'h37b7;
aud[20007]=16'h37c2;
aud[20008]=16'h37cc;
aud[20009]=16'h37d7;
aud[20010]=16'h37e1;
aud[20011]=16'h37ec;
aud[20012]=16'h37f6;
aud[20013]=16'h3801;
aud[20014]=16'h380b;
aud[20015]=16'h3815;
aud[20016]=16'h3820;
aud[20017]=16'h382a;
aud[20018]=16'h3834;
aud[20019]=16'h383f;
aud[20020]=16'h3849;
aud[20021]=16'h3853;
aud[20022]=16'h385d;
aud[20023]=16'h3867;
aud[20024]=16'h3871;
aud[20025]=16'h387b;
aud[20026]=16'h3886;
aud[20027]=16'h3890;
aud[20028]=16'h389a;
aud[20029]=16'h38a4;
aud[20030]=16'h38ae;
aud[20031]=16'h38b8;
aud[20032]=16'h38c1;
aud[20033]=16'h38cb;
aud[20034]=16'h38d5;
aud[20035]=16'h38df;
aud[20036]=16'h38e9;
aud[20037]=16'h38f3;
aud[20038]=16'h38fd;
aud[20039]=16'h3906;
aud[20040]=16'h3910;
aud[20041]=16'h391a;
aud[20042]=16'h3923;
aud[20043]=16'h392d;
aud[20044]=16'h3937;
aud[20045]=16'h3940;
aud[20046]=16'h394a;
aud[20047]=16'h3953;
aud[20048]=16'h395d;
aud[20049]=16'h3966;
aud[20050]=16'h3970;
aud[20051]=16'h3979;
aud[20052]=16'h3983;
aud[20053]=16'h398c;
aud[20054]=16'h3995;
aud[20055]=16'h399f;
aud[20056]=16'h39a8;
aud[20057]=16'h39b1;
aud[20058]=16'h39bb;
aud[20059]=16'h39c4;
aud[20060]=16'h39cd;
aud[20061]=16'h39d6;
aud[20062]=16'h39e0;
aud[20063]=16'h39e9;
aud[20064]=16'h39f2;
aud[20065]=16'h39fb;
aud[20066]=16'h3a04;
aud[20067]=16'h3a0d;
aud[20068]=16'h3a16;
aud[20069]=16'h3a1f;
aud[20070]=16'h3a28;
aud[20071]=16'h3a31;
aud[20072]=16'h3a3a;
aud[20073]=16'h3a43;
aud[20074]=16'h3a4c;
aud[20075]=16'h3a54;
aud[20076]=16'h3a5d;
aud[20077]=16'h3a66;
aud[20078]=16'h3a6f;
aud[20079]=16'h3a78;
aud[20080]=16'h3a80;
aud[20081]=16'h3a89;
aud[20082]=16'h3a92;
aud[20083]=16'h3a9a;
aud[20084]=16'h3aa3;
aud[20085]=16'h3aab;
aud[20086]=16'h3ab4;
aud[20087]=16'h3abc;
aud[20088]=16'h3ac5;
aud[20089]=16'h3acd;
aud[20090]=16'h3ad6;
aud[20091]=16'h3ade;
aud[20092]=16'h3ae7;
aud[20093]=16'h3aef;
aud[20094]=16'h3af7;
aud[20095]=16'h3b00;
aud[20096]=16'h3b08;
aud[20097]=16'h3b10;
aud[20098]=16'h3b19;
aud[20099]=16'h3b21;
aud[20100]=16'h3b29;
aud[20101]=16'h3b31;
aud[20102]=16'h3b39;
aud[20103]=16'h3b41;
aud[20104]=16'h3b4a;
aud[20105]=16'h3b52;
aud[20106]=16'h3b5a;
aud[20107]=16'h3b62;
aud[20108]=16'h3b6a;
aud[20109]=16'h3b72;
aud[20110]=16'h3b7a;
aud[20111]=16'h3b81;
aud[20112]=16'h3b89;
aud[20113]=16'h3b91;
aud[20114]=16'h3b99;
aud[20115]=16'h3ba1;
aud[20116]=16'h3ba9;
aud[20117]=16'h3bb0;
aud[20118]=16'h3bb8;
aud[20119]=16'h3bc0;
aud[20120]=16'h3bc7;
aud[20121]=16'h3bcf;
aud[20122]=16'h3bd7;
aud[20123]=16'h3bde;
aud[20124]=16'h3be6;
aud[20125]=16'h3bed;
aud[20126]=16'h3bf5;
aud[20127]=16'h3bfc;
aud[20128]=16'h3c04;
aud[20129]=16'h3c0b;
aud[20130]=16'h3c13;
aud[20131]=16'h3c1a;
aud[20132]=16'h3c21;
aud[20133]=16'h3c29;
aud[20134]=16'h3c30;
aud[20135]=16'h3c37;
aud[20136]=16'h3c3f;
aud[20137]=16'h3c46;
aud[20138]=16'h3c4d;
aud[20139]=16'h3c54;
aud[20140]=16'h3c5b;
aud[20141]=16'h3c63;
aud[20142]=16'h3c6a;
aud[20143]=16'h3c71;
aud[20144]=16'h3c78;
aud[20145]=16'h3c7f;
aud[20146]=16'h3c86;
aud[20147]=16'h3c8d;
aud[20148]=16'h3c94;
aud[20149]=16'h3c9b;
aud[20150]=16'h3ca1;
aud[20151]=16'h3ca8;
aud[20152]=16'h3caf;
aud[20153]=16'h3cb6;
aud[20154]=16'h3cbd;
aud[20155]=16'h3cc3;
aud[20156]=16'h3cca;
aud[20157]=16'h3cd1;
aud[20158]=16'h3cd7;
aud[20159]=16'h3cde;
aud[20160]=16'h3ce5;
aud[20161]=16'h3ceb;
aud[20162]=16'h3cf2;
aud[20163]=16'h3cf8;
aud[20164]=16'h3cff;
aud[20165]=16'h3d05;
aud[20166]=16'h3d0c;
aud[20167]=16'h3d12;
aud[20168]=16'h3d19;
aud[20169]=16'h3d1f;
aud[20170]=16'h3d25;
aud[20171]=16'h3d2c;
aud[20172]=16'h3d32;
aud[20173]=16'h3d38;
aud[20174]=16'h3d3f;
aud[20175]=16'h3d45;
aud[20176]=16'h3d4b;
aud[20177]=16'h3d51;
aud[20178]=16'h3d57;
aud[20179]=16'h3d5d;
aud[20180]=16'h3d63;
aud[20181]=16'h3d69;
aud[20182]=16'h3d6f;
aud[20183]=16'h3d75;
aud[20184]=16'h3d7b;
aud[20185]=16'h3d81;
aud[20186]=16'h3d87;
aud[20187]=16'h3d8d;
aud[20188]=16'h3d93;
aud[20189]=16'h3d99;
aud[20190]=16'h3d9f;
aud[20191]=16'h3da4;
aud[20192]=16'h3daa;
aud[20193]=16'h3db0;
aud[20194]=16'h3db6;
aud[20195]=16'h3dbb;
aud[20196]=16'h3dc1;
aud[20197]=16'h3dc7;
aud[20198]=16'h3dcc;
aud[20199]=16'h3dd2;
aud[20200]=16'h3dd7;
aud[20201]=16'h3ddd;
aud[20202]=16'h3de2;
aud[20203]=16'h3de8;
aud[20204]=16'h3ded;
aud[20205]=16'h3df3;
aud[20206]=16'h3df8;
aud[20207]=16'h3dfd;
aud[20208]=16'h3e03;
aud[20209]=16'h3e08;
aud[20210]=16'h3e0d;
aud[20211]=16'h3e12;
aud[20212]=16'h3e18;
aud[20213]=16'h3e1d;
aud[20214]=16'h3e22;
aud[20215]=16'h3e27;
aud[20216]=16'h3e2c;
aud[20217]=16'h3e31;
aud[20218]=16'h3e36;
aud[20219]=16'h3e3b;
aud[20220]=16'h3e40;
aud[20221]=16'h3e45;
aud[20222]=16'h3e4a;
aud[20223]=16'h3e4f;
aud[20224]=16'h3e54;
aud[20225]=16'h3e59;
aud[20226]=16'h3e5e;
aud[20227]=16'h3e62;
aud[20228]=16'h3e67;
aud[20229]=16'h3e6c;
aud[20230]=16'h3e71;
aud[20231]=16'h3e75;
aud[20232]=16'h3e7a;
aud[20233]=16'h3e7f;
aud[20234]=16'h3e83;
aud[20235]=16'h3e88;
aud[20236]=16'h3e8c;
aud[20237]=16'h3e91;
aud[20238]=16'h3e95;
aud[20239]=16'h3e9a;
aud[20240]=16'h3e9e;
aud[20241]=16'h3ea3;
aud[20242]=16'h3ea7;
aud[20243]=16'h3eac;
aud[20244]=16'h3eb0;
aud[20245]=16'h3eb4;
aud[20246]=16'h3eb9;
aud[20247]=16'h3ebd;
aud[20248]=16'h3ec1;
aud[20249]=16'h3ec5;
aud[20250]=16'h3ec9;
aud[20251]=16'h3ecd;
aud[20252]=16'h3ed2;
aud[20253]=16'h3ed6;
aud[20254]=16'h3eda;
aud[20255]=16'h3ede;
aud[20256]=16'h3ee2;
aud[20257]=16'h3ee6;
aud[20258]=16'h3eea;
aud[20259]=16'h3eee;
aud[20260]=16'h3ef2;
aud[20261]=16'h3ef5;
aud[20262]=16'h3ef9;
aud[20263]=16'h3efd;
aud[20264]=16'h3f01;
aud[20265]=16'h3f05;
aud[20266]=16'h3f08;
aud[20267]=16'h3f0c;
aud[20268]=16'h3f10;
aud[20269]=16'h3f13;
aud[20270]=16'h3f17;
aud[20271]=16'h3f1b;
aud[20272]=16'h3f1e;
aud[20273]=16'h3f22;
aud[20274]=16'h3f25;
aud[20275]=16'h3f29;
aud[20276]=16'h3f2c;
aud[20277]=16'h3f30;
aud[20278]=16'h3f33;
aud[20279]=16'h3f36;
aud[20280]=16'h3f3a;
aud[20281]=16'h3f3d;
aud[20282]=16'h3f40;
aud[20283]=16'h3f43;
aud[20284]=16'h3f47;
aud[20285]=16'h3f4a;
aud[20286]=16'h3f4d;
aud[20287]=16'h3f50;
aud[20288]=16'h3f53;
aud[20289]=16'h3f56;
aud[20290]=16'h3f5a;
aud[20291]=16'h3f5d;
aud[20292]=16'h3f60;
aud[20293]=16'h3f63;
aud[20294]=16'h3f65;
aud[20295]=16'h3f68;
aud[20296]=16'h3f6b;
aud[20297]=16'h3f6e;
aud[20298]=16'h3f71;
aud[20299]=16'h3f74;
aud[20300]=16'h3f77;
aud[20301]=16'h3f79;
aud[20302]=16'h3f7c;
aud[20303]=16'h3f7f;
aud[20304]=16'h3f81;
aud[20305]=16'h3f84;
aud[20306]=16'h3f87;
aud[20307]=16'h3f89;
aud[20308]=16'h3f8c;
aud[20309]=16'h3f8e;
aud[20310]=16'h3f91;
aud[20311]=16'h3f93;
aud[20312]=16'h3f96;
aud[20313]=16'h3f98;
aud[20314]=16'h3f9b;
aud[20315]=16'h3f9d;
aud[20316]=16'h3f9f;
aud[20317]=16'h3fa2;
aud[20318]=16'h3fa4;
aud[20319]=16'h3fa6;
aud[20320]=16'h3fa8;
aud[20321]=16'h3fab;
aud[20322]=16'h3fad;
aud[20323]=16'h3faf;
aud[20324]=16'h3fb1;
aud[20325]=16'h3fb3;
aud[20326]=16'h3fb5;
aud[20327]=16'h3fb7;
aud[20328]=16'h3fb9;
aud[20329]=16'h3fbb;
aud[20330]=16'h3fbd;
aud[20331]=16'h3fbf;
aud[20332]=16'h3fc1;
aud[20333]=16'h3fc3;
aud[20334]=16'h3fc5;
aud[20335]=16'h3fc7;
aud[20336]=16'h3fc8;
aud[20337]=16'h3fca;
aud[20338]=16'h3fcc;
aud[20339]=16'h3fcd;
aud[20340]=16'h3fcf;
aud[20341]=16'h3fd1;
aud[20342]=16'h3fd2;
aud[20343]=16'h3fd4;
aud[20344]=16'h3fd6;
aud[20345]=16'h3fd7;
aud[20346]=16'h3fd9;
aud[20347]=16'h3fda;
aud[20348]=16'h3fdc;
aud[20349]=16'h3fdd;
aud[20350]=16'h3fde;
aud[20351]=16'h3fe0;
aud[20352]=16'h3fe1;
aud[20353]=16'h3fe2;
aud[20354]=16'h3fe4;
aud[20355]=16'h3fe5;
aud[20356]=16'h3fe6;
aud[20357]=16'h3fe7;
aud[20358]=16'h3fe8;
aud[20359]=16'h3fea;
aud[20360]=16'h3feb;
aud[20361]=16'h3fec;
aud[20362]=16'h3fed;
aud[20363]=16'h3fee;
aud[20364]=16'h3fef;
aud[20365]=16'h3ff0;
aud[20366]=16'h3ff1;
aud[20367]=16'h3ff2;
aud[20368]=16'h3ff3;
aud[20369]=16'h3ff3;
aud[20370]=16'h3ff4;
aud[20371]=16'h3ff5;
aud[20372]=16'h3ff6;
aud[20373]=16'h3ff7;
aud[20374]=16'h3ff7;
aud[20375]=16'h3ff8;
aud[20376]=16'h3ff9;
aud[20377]=16'h3ff9;
aud[20378]=16'h3ffa;
aud[20379]=16'h3ffa;
aud[20380]=16'h3ffb;
aud[20381]=16'h3ffb;
aud[20382]=16'h3ffc;
aud[20383]=16'h3ffc;
aud[20384]=16'h3ffd;
aud[20385]=16'h3ffd;
aud[20386]=16'h3ffe;
aud[20387]=16'h3ffe;
aud[20388]=16'h3ffe;
aud[20389]=16'h3fff;
aud[20390]=16'h3fff;
aud[20391]=16'h3fff;
aud[20392]=16'h3fff;
aud[20393]=16'h3fff;
aud[20394]=16'h4000;
aud[20395]=16'h4000;
aud[20396]=16'h4000;
aud[20397]=16'h4000;
aud[20398]=16'h4000;
aud[20399]=16'h4000;
aud[20400]=16'h4000;
aud[20401]=16'h4000;
aud[20402]=16'h4000;
aud[20403]=16'h4000;
aud[20404]=16'h4000;
aud[20405]=16'h3fff;
aud[20406]=16'h3fff;
aud[20407]=16'h3fff;
aud[20408]=16'h3fff;
aud[20409]=16'h3fff;
aud[20410]=16'h3ffe;
aud[20411]=16'h3ffe;
aud[20412]=16'h3ffe;
aud[20413]=16'h3ffd;
aud[20414]=16'h3ffd;
aud[20415]=16'h3ffc;
aud[20416]=16'h3ffc;
aud[20417]=16'h3ffb;
aud[20418]=16'h3ffb;
aud[20419]=16'h3ffa;
aud[20420]=16'h3ffa;
aud[20421]=16'h3ff9;
aud[20422]=16'h3ff9;
aud[20423]=16'h3ff8;
aud[20424]=16'h3ff7;
aud[20425]=16'h3ff7;
aud[20426]=16'h3ff6;
aud[20427]=16'h3ff5;
aud[20428]=16'h3ff4;
aud[20429]=16'h3ff3;
aud[20430]=16'h3ff3;
aud[20431]=16'h3ff2;
aud[20432]=16'h3ff1;
aud[20433]=16'h3ff0;
aud[20434]=16'h3fef;
aud[20435]=16'h3fee;
aud[20436]=16'h3fed;
aud[20437]=16'h3fec;
aud[20438]=16'h3feb;
aud[20439]=16'h3fea;
aud[20440]=16'h3fe8;
aud[20441]=16'h3fe7;
aud[20442]=16'h3fe6;
aud[20443]=16'h3fe5;
aud[20444]=16'h3fe4;
aud[20445]=16'h3fe2;
aud[20446]=16'h3fe1;
aud[20447]=16'h3fe0;
aud[20448]=16'h3fde;
aud[20449]=16'h3fdd;
aud[20450]=16'h3fdc;
aud[20451]=16'h3fda;
aud[20452]=16'h3fd9;
aud[20453]=16'h3fd7;
aud[20454]=16'h3fd6;
aud[20455]=16'h3fd4;
aud[20456]=16'h3fd2;
aud[20457]=16'h3fd1;
aud[20458]=16'h3fcf;
aud[20459]=16'h3fcd;
aud[20460]=16'h3fcc;
aud[20461]=16'h3fca;
aud[20462]=16'h3fc8;
aud[20463]=16'h3fc7;
aud[20464]=16'h3fc5;
aud[20465]=16'h3fc3;
aud[20466]=16'h3fc1;
aud[20467]=16'h3fbf;
aud[20468]=16'h3fbd;
aud[20469]=16'h3fbb;
aud[20470]=16'h3fb9;
aud[20471]=16'h3fb7;
aud[20472]=16'h3fb5;
aud[20473]=16'h3fb3;
aud[20474]=16'h3fb1;
aud[20475]=16'h3faf;
aud[20476]=16'h3fad;
aud[20477]=16'h3fab;
aud[20478]=16'h3fa8;
aud[20479]=16'h3fa6;
aud[20480]=16'h3fa4;
aud[20481]=16'h3fa2;
aud[20482]=16'h3f9f;
aud[20483]=16'h3f9d;
aud[20484]=16'h3f9b;
aud[20485]=16'h3f98;
aud[20486]=16'h3f96;
aud[20487]=16'h3f93;
aud[20488]=16'h3f91;
aud[20489]=16'h3f8e;
aud[20490]=16'h3f8c;
aud[20491]=16'h3f89;
aud[20492]=16'h3f87;
aud[20493]=16'h3f84;
aud[20494]=16'h3f81;
aud[20495]=16'h3f7f;
aud[20496]=16'h3f7c;
aud[20497]=16'h3f79;
aud[20498]=16'h3f77;
aud[20499]=16'h3f74;
aud[20500]=16'h3f71;
aud[20501]=16'h3f6e;
aud[20502]=16'h3f6b;
aud[20503]=16'h3f68;
aud[20504]=16'h3f65;
aud[20505]=16'h3f63;
aud[20506]=16'h3f60;
aud[20507]=16'h3f5d;
aud[20508]=16'h3f5a;
aud[20509]=16'h3f56;
aud[20510]=16'h3f53;
aud[20511]=16'h3f50;
aud[20512]=16'h3f4d;
aud[20513]=16'h3f4a;
aud[20514]=16'h3f47;
aud[20515]=16'h3f43;
aud[20516]=16'h3f40;
aud[20517]=16'h3f3d;
aud[20518]=16'h3f3a;
aud[20519]=16'h3f36;
aud[20520]=16'h3f33;
aud[20521]=16'h3f30;
aud[20522]=16'h3f2c;
aud[20523]=16'h3f29;
aud[20524]=16'h3f25;
aud[20525]=16'h3f22;
aud[20526]=16'h3f1e;
aud[20527]=16'h3f1b;
aud[20528]=16'h3f17;
aud[20529]=16'h3f13;
aud[20530]=16'h3f10;
aud[20531]=16'h3f0c;
aud[20532]=16'h3f08;
aud[20533]=16'h3f05;
aud[20534]=16'h3f01;
aud[20535]=16'h3efd;
aud[20536]=16'h3ef9;
aud[20537]=16'h3ef5;
aud[20538]=16'h3ef2;
aud[20539]=16'h3eee;
aud[20540]=16'h3eea;
aud[20541]=16'h3ee6;
aud[20542]=16'h3ee2;
aud[20543]=16'h3ede;
aud[20544]=16'h3eda;
aud[20545]=16'h3ed6;
aud[20546]=16'h3ed2;
aud[20547]=16'h3ecd;
aud[20548]=16'h3ec9;
aud[20549]=16'h3ec5;
aud[20550]=16'h3ec1;
aud[20551]=16'h3ebd;
aud[20552]=16'h3eb9;
aud[20553]=16'h3eb4;
aud[20554]=16'h3eb0;
aud[20555]=16'h3eac;
aud[20556]=16'h3ea7;
aud[20557]=16'h3ea3;
aud[20558]=16'h3e9e;
aud[20559]=16'h3e9a;
aud[20560]=16'h3e95;
aud[20561]=16'h3e91;
aud[20562]=16'h3e8c;
aud[20563]=16'h3e88;
aud[20564]=16'h3e83;
aud[20565]=16'h3e7f;
aud[20566]=16'h3e7a;
aud[20567]=16'h3e75;
aud[20568]=16'h3e71;
aud[20569]=16'h3e6c;
aud[20570]=16'h3e67;
aud[20571]=16'h3e62;
aud[20572]=16'h3e5e;
aud[20573]=16'h3e59;
aud[20574]=16'h3e54;
aud[20575]=16'h3e4f;
aud[20576]=16'h3e4a;
aud[20577]=16'h3e45;
aud[20578]=16'h3e40;
aud[20579]=16'h3e3b;
aud[20580]=16'h3e36;
aud[20581]=16'h3e31;
aud[20582]=16'h3e2c;
aud[20583]=16'h3e27;
aud[20584]=16'h3e22;
aud[20585]=16'h3e1d;
aud[20586]=16'h3e18;
aud[20587]=16'h3e12;
aud[20588]=16'h3e0d;
aud[20589]=16'h3e08;
aud[20590]=16'h3e03;
aud[20591]=16'h3dfd;
aud[20592]=16'h3df8;
aud[20593]=16'h3df3;
aud[20594]=16'h3ded;
aud[20595]=16'h3de8;
aud[20596]=16'h3de2;
aud[20597]=16'h3ddd;
aud[20598]=16'h3dd7;
aud[20599]=16'h3dd2;
aud[20600]=16'h3dcc;
aud[20601]=16'h3dc7;
aud[20602]=16'h3dc1;
aud[20603]=16'h3dbb;
aud[20604]=16'h3db6;
aud[20605]=16'h3db0;
aud[20606]=16'h3daa;
aud[20607]=16'h3da4;
aud[20608]=16'h3d9f;
aud[20609]=16'h3d99;
aud[20610]=16'h3d93;
aud[20611]=16'h3d8d;
aud[20612]=16'h3d87;
aud[20613]=16'h3d81;
aud[20614]=16'h3d7b;
aud[20615]=16'h3d75;
aud[20616]=16'h3d6f;
aud[20617]=16'h3d69;
aud[20618]=16'h3d63;
aud[20619]=16'h3d5d;
aud[20620]=16'h3d57;
aud[20621]=16'h3d51;
aud[20622]=16'h3d4b;
aud[20623]=16'h3d45;
aud[20624]=16'h3d3f;
aud[20625]=16'h3d38;
aud[20626]=16'h3d32;
aud[20627]=16'h3d2c;
aud[20628]=16'h3d25;
aud[20629]=16'h3d1f;
aud[20630]=16'h3d19;
aud[20631]=16'h3d12;
aud[20632]=16'h3d0c;
aud[20633]=16'h3d05;
aud[20634]=16'h3cff;
aud[20635]=16'h3cf8;
aud[20636]=16'h3cf2;
aud[20637]=16'h3ceb;
aud[20638]=16'h3ce5;
aud[20639]=16'h3cde;
aud[20640]=16'h3cd7;
aud[20641]=16'h3cd1;
aud[20642]=16'h3cca;
aud[20643]=16'h3cc3;
aud[20644]=16'h3cbd;
aud[20645]=16'h3cb6;
aud[20646]=16'h3caf;
aud[20647]=16'h3ca8;
aud[20648]=16'h3ca1;
aud[20649]=16'h3c9b;
aud[20650]=16'h3c94;
aud[20651]=16'h3c8d;
aud[20652]=16'h3c86;
aud[20653]=16'h3c7f;
aud[20654]=16'h3c78;
aud[20655]=16'h3c71;
aud[20656]=16'h3c6a;
aud[20657]=16'h3c63;
aud[20658]=16'h3c5b;
aud[20659]=16'h3c54;
aud[20660]=16'h3c4d;
aud[20661]=16'h3c46;
aud[20662]=16'h3c3f;
aud[20663]=16'h3c37;
aud[20664]=16'h3c30;
aud[20665]=16'h3c29;
aud[20666]=16'h3c21;
aud[20667]=16'h3c1a;
aud[20668]=16'h3c13;
aud[20669]=16'h3c0b;
aud[20670]=16'h3c04;
aud[20671]=16'h3bfc;
aud[20672]=16'h3bf5;
aud[20673]=16'h3bed;
aud[20674]=16'h3be6;
aud[20675]=16'h3bde;
aud[20676]=16'h3bd7;
aud[20677]=16'h3bcf;
aud[20678]=16'h3bc7;
aud[20679]=16'h3bc0;
aud[20680]=16'h3bb8;
aud[20681]=16'h3bb0;
aud[20682]=16'h3ba9;
aud[20683]=16'h3ba1;
aud[20684]=16'h3b99;
aud[20685]=16'h3b91;
aud[20686]=16'h3b89;
aud[20687]=16'h3b81;
aud[20688]=16'h3b7a;
aud[20689]=16'h3b72;
aud[20690]=16'h3b6a;
aud[20691]=16'h3b62;
aud[20692]=16'h3b5a;
aud[20693]=16'h3b52;
aud[20694]=16'h3b4a;
aud[20695]=16'h3b41;
aud[20696]=16'h3b39;
aud[20697]=16'h3b31;
aud[20698]=16'h3b29;
aud[20699]=16'h3b21;
aud[20700]=16'h3b19;
aud[20701]=16'h3b10;
aud[20702]=16'h3b08;
aud[20703]=16'h3b00;
aud[20704]=16'h3af7;
aud[20705]=16'h3aef;
aud[20706]=16'h3ae7;
aud[20707]=16'h3ade;
aud[20708]=16'h3ad6;
aud[20709]=16'h3acd;
aud[20710]=16'h3ac5;
aud[20711]=16'h3abc;
aud[20712]=16'h3ab4;
aud[20713]=16'h3aab;
aud[20714]=16'h3aa3;
aud[20715]=16'h3a9a;
aud[20716]=16'h3a92;
aud[20717]=16'h3a89;
aud[20718]=16'h3a80;
aud[20719]=16'h3a78;
aud[20720]=16'h3a6f;
aud[20721]=16'h3a66;
aud[20722]=16'h3a5d;
aud[20723]=16'h3a54;
aud[20724]=16'h3a4c;
aud[20725]=16'h3a43;
aud[20726]=16'h3a3a;
aud[20727]=16'h3a31;
aud[20728]=16'h3a28;
aud[20729]=16'h3a1f;
aud[20730]=16'h3a16;
aud[20731]=16'h3a0d;
aud[20732]=16'h3a04;
aud[20733]=16'h39fb;
aud[20734]=16'h39f2;
aud[20735]=16'h39e9;
aud[20736]=16'h39e0;
aud[20737]=16'h39d6;
aud[20738]=16'h39cd;
aud[20739]=16'h39c4;
aud[20740]=16'h39bb;
aud[20741]=16'h39b1;
aud[20742]=16'h39a8;
aud[20743]=16'h399f;
aud[20744]=16'h3995;
aud[20745]=16'h398c;
aud[20746]=16'h3983;
aud[20747]=16'h3979;
aud[20748]=16'h3970;
aud[20749]=16'h3966;
aud[20750]=16'h395d;
aud[20751]=16'h3953;
aud[20752]=16'h394a;
aud[20753]=16'h3940;
aud[20754]=16'h3937;
aud[20755]=16'h392d;
aud[20756]=16'h3923;
aud[20757]=16'h391a;
aud[20758]=16'h3910;
aud[20759]=16'h3906;
aud[20760]=16'h38fd;
aud[20761]=16'h38f3;
aud[20762]=16'h38e9;
aud[20763]=16'h38df;
aud[20764]=16'h38d5;
aud[20765]=16'h38cb;
aud[20766]=16'h38c1;
aud[20767]=16'h38b8;
aud[20768]=16'h38ae;
aud[20769]=16'h38a4;
aud[20770]=16'h389a;
aud[20771]=16'h3890;
aud[20772]=16'h3886;
aud[20773]=16'h387b;
aud[20774]=16'h3871;
aud[20775]=16'h3867;
aud[20776]=16'h385d;
aud[20777]=16'h3853;
aud[20778]=16'h3849;
aud[20779]=16'h383f;
aud[20780]=16'h3834;
aud[20781]=16'h382a;
aud[20782]=16'h3820;
aud[20783]=16'h3815;
aud[20784]=16'h380b;
aud[20785]=16'h3801;
aud[20786]=16'h37f6;
aud[20787]=16'h37ec;
aud[20788]=16'h37e1;
aud[20789]=16'h37d7;
aud[20790]=16'h37cc;
aud[20791]=16'h37c2;
aud[20792]=16'h37b7;
aud[20793]=16'h37ad;
aud[20794]=16'h37a2;
aud[20795]=16'h3798;
aud[20796]=16'h378d;
aud[20797]=16'h3782;
aud[20798]=16'h3778;
aud[20799]=16'h376d;
aud[20800]=16'h3762;
aud[20801]=16'h3757;
aud[20802]=16'h374d;
aud[20803]=16'h3742;
aud[20804]=16'h3737;
aud[20805]=16'h372c;
aud[20806]=16'h3721;
aud[20807]=16'h3716;
aud[20808]=16'h370b;
aud[20809]=16'h3701;
aud[20810]=16'h36f6;
aud[20811]=16'h36eb;
aud[20812]=16'h36e0;
aud[20813]=16'h36d4;
aud[20814]=16'h36c9;
aud[20815]=16'h36be;
aud[20816]=16'h36b3;
aud[20817]=16'h36a8;
aud[20818]=16'h369d;
aud[20819]=16'h3692;
aud[20820]=16'h3686;
aud[20821]=16'h367b;
aud[20822]=16'h3670;
aud[20823]=16'h3665;
aud[20824]=16'h3659;
aud[20825]=16'h364e;
aud[20826]=16'h3643;
aud[20827]=16'h3637;
aud[20828]=16'h362c;
aud[20829]=16'h3620;
aud[20830]=16'h3615;
aud[20831]=16'h3609;
aud[20832]=16'h35fe;
aud[20833]=16'h35f2;
aud[20834]=16'h35e7;
aud[20835]=16'h35db;
aud[20836]=16'h35d0;
aud[20837]=16'h35c4;
aud[20838]=16'h35b8;
aud[20839]=16'h35ad;
aud[20840]=16'h35a1;
aud[20841]=16'h3595;
aud[20842]=16'h358a;
aud[20843]=16'h357e;
aud[20844]=16'h3572;
aud[20845]=16'h3566;
aud[20846]=16'h355a;
aud[20847]=16'h354f;
aud[20848]=16'h3543;
aud[20849]=16'h3537;
aud[20850]=16'h352b;
aud[20851]=16'h351f;
aud[20852]=16'h3513;
aud[20853]=16'h3507;
aud[20854]=16'h34fb;
aud[20855]=16'h34ef;
aud[20856]=16'h34e3;
aud[20857]=16'h34d7;
aud[20858]=16'h34cb;
aud[20859]=16'h34be;
aud[20860]=16'h34b2;
aud[20861]=16'h34a6;
aud[20862]=16'h349a;
aud[20863]=16'h348e;
aud[20864]=16'h3481;
aud[20865]=16'h3475;
aud[20866]=16'h3469;
aud[20867]=16'h345d;
aud[20868]=16'h3450;
aud[20869]=16'h3444;
aud[20870]=16'h3437;
aud[20871]=16'h342b;
aud[20872]=16'h341f;
aud[20873]=16'h3412;
aud[20874]=16'h3406;
aud[20875]=16'h33f9;
aud[20876]=16'h33ed;
aud[20877]=16'h33e0;
aud[20878]=16'h33d4;
aud[20879]=16'h33c7;
aud[20880]=16'h33ba;
aud[20881]=16'h33ae;
aud[20882]=16'h33a1;
aud[20883]=16'h3394;
aud[20884]=16'h3388;
aud[20885]=16'h337b;
aud[20886]=16'h336e;
aud[20887]=16'h3361;
aud[20888]=16'h3355;
aud[20889]=16'h3348;
aud[20890]=16'h333b;
aud[20891]=16'h332e;
aud[20892]=16'h3321;
aud[20893]=16'h3314;
aud[20894]=16'h3307;
aud[20895]=16'h32fa;
aud[20896]=16'h32ed;
aud[20897]=16'h32e0;
aud[20898]=16'h32d3;
aud[20899]=16'h32c6;
aud[20900]=16'h32b9;
aud[20901]=16'h32ac;
aud[20902]=16'h329f;
aud[20903]=16'h3292;
aud[20904]=16'h3285;
aud[20905]=16'h3278;
aud[20906]=16'h326a;
aud[20907]=16'h325d;
aud[20908]=16'h3250;
aud[20909]=16'h3243;
aud[20910]=16'h3235;
aud[20911]=16'h3228;
aud[20912]=16'h321b;
aud[20913]=16'h320d;
aud[20914]=16'h3200;
aud[20915]=16'h31f3;
aud[20916]=16'h31e5;
aud[20917]=16'h31d8;
aud[20918]=16'h31ca;
aud[20919]=16'h31bd;
aud[20920]=16'h31af;
aud[20921]=16'h31a2;
aud[20922]=16'h3194;
aud[20923]=16'h3187;
aud[20924]=16'h3179;
aud[20925]=16'h316b;
aud[20926]=16'h315e;
aud[20927]=16'h3150;
aud[20928]=16'h3142;
aud[20929]=16'h3135;
aud[20930]=16'h3127;
aud[20931]=16'h3119;
aud[20932]=16'h310b;
aud[20933]=16'h30fe;
aud[20934]=16'h30f0;
aud[20935]=16'h30e2;
aud[20936]=16'h30d4;
aud[20937]=16'h30c6;
aud[20938]=16'h30b8;
aud[20939]=16'h30aa;
aud[20940]=16'h309d;
aud[20941]=16'h308f;
aud[20942]=16'h3081;
aud[20943]=16'h3073;
aud[20944]=16'h3065;
aud[20945]=16'h3057;
aud[20946]=16'h3048;
aud[20947]=16'h303a;
aud[20948]=16'h302c;
aud[20949]=16'h301e;
aud[20950]=16'h3010;
aud[20951]=16'h3002;
aud[20952]=16'h2ff4;
aud[20953]=16'h2fe5;
aud[20954]=16'h2fd7;
aud[20955]=16'h2fc9;
aud[20956]=16'h2fbb;
aud[20957]=16'h2fac;
aud[20958]=16'h2f9e;
aud[20959]=16'h2f90;
aud[20960]=16'h2f81;
aud[20961]=16'h2f73;
aud[20962]=16'h2f65;
aud[20963]=16'h2f56;
aud[20964]=16'h2f48;
aud[20965]=16'h2f39;
aud[20966]=16'h2f2b;
aud[20967]=16'h2f1c;
aud[20968]=16'h2f0e;
aud[20969]=16'h2eff;
aud[20970]=16'h2ef1;
aud[20971]=16'h2ee2;
aud[20972]=16'h2ed3;
aud[20973]=16'h2ec5;
aud[20974]=16'h2eb6;
aud[20975]=16'h2ea7;
aud[20976]=16'h2e99;
aud[20977]=16'h2e8a;
aud[20978]=16'h2e7b;
aud[20979]=16'h2e6d;
aud[20980]=16'h2e5e;
aud[20981]=16'h2e4f;
aud[20982]=16'h2e40;
aud[20983]=16'h2e31;
aud[20984]=16'h2e22;
aud[20985]=16'h2e14;
aud[20986]=16'h2e05;
aud[20987]=16'h2df6;
aud[20988]=16'h2de7;
aud[20989]=16'h2dd8;
aud[20990]=16'h2dc9;
aud[20991]=16'h2dba;
aud[20992]=16'h2dab;
aud[20993]=16'h2d9c;
aud[20994]=16'h2d8d;
aud[20995]=16'h2d7e;
aud[20996]=16'h2d6f;
aud[20997]=16'h2d60;
aud[20998]=16'h2d50;
aud[20999]=16'h2d41;
aud[21000]=16'h2d32;
aud[21001]=16'h2d23;
aud[21002]=16'h2d14;
aud[21003]=16'h2d04;
aud[21004]=16'h2cf5;
aud[21005]=16'h2ce6;
aud[21006]=16'h2cd7;
aud[21007]=16'h2cc7;
aud[21008]=16'h2cb8;
aud[21009]=16'h2ca9;
aud[21010]=16'h2c99;
aud[21011]=16'h2c8a;
aud[21012]=16'h2c7a;
aud[21013]=16'h2c6b;
aud[21014]=16'h2c5c;
aud[21015]=16'h2c4c;
aud[21016]=16'h2c3d;
aud[21017]=16'h2c2d;
aud[21018]=16'h2c1e;
aud[21019]=16'h2c0e;
aud[21020]=16'h2bfe;
aud[21021]=16'h2bef;
aud[21022]=16'h2bdf;
aud[21023]=16'h2bd0;
aud[21024]=16'h2bc0;
aud[21025]=16'h2bb0;
aud[21026]=16'h2ba1;
aud[21027]=16'h2b91;
aud[21028]=16'h2b81;
aud[21029]=16'h2b71;
aud[21030]=16'h2b62;
aud[21031]=16'h2b52;
aud[21032]=16'h2b42;
aud[21033]=16'h2b32;
aud[21034]=16'h2b22;
aud[21035]=16'h2b13;
aud[21036]=16'h2b03;
aud[21037]=16'h2af3;
aud[21038]=16'h2ae3;
aud[21039]=16'h2ad3;
aud[21040]=16'h2ac3;
aud[21041]=16'h2ab3;
aud[21042]=16'h2aa3;
aud[21043]=16'h2a93;
aud[21044]=16'h2a83;
aud[21045]=16'h2a73;
aud[21046]=16'h2a63;
aud[21047]=16'h2a53;
aud[21048]=16'h2a43;
aud[21049]=16'h2a33;
aud[21050]=16'h2a23;
aud[21051]=16'h2a12;
aud[21052]=16'h2a02;
aud[21053]=16'h29f2;
aud[21054]=16'h29e2;
aud[21055]=16'h29d2;
aud[21056]=16'h29c1;
aud[21057]=16'h29b1;
aud[21058]=16'h29a1;
aud[21059]=16'h2991;
aud[21060]=16'h2980;
aud[21061]=16'h2970;
aud[21062]=16'h2960;
aud[21063]=16'h294f;
aud[21064]=16'h293f;
aud[21065]=16'h292e;
aud[21066]=16'h291e;
aud[21067]=16'h290e;
aud[21068]=16'h28fd;
aud[21069]=16'h28ed;
aud[21070]=16'h28dc;
aud[21071]=16'h28cc;
aud[21072]=16'h28bb;
aud[21073]=16'h28aa;
aud[21074]=16'h289a;
aud[21075]=16'h2889;
aud[21076]=16'h2879;
aud[21077]=16'h2868;
aud[21078]=16'h2857;
aud[21079]=16'h2847;
aud[21080]=16'h2836;
aud[21081]=16'h2825;
aud[21082]=16'h2815;
aud[21083]=16'h2804;
aud[21084]=16'h27f3;
aud[21085]=16'h27e2;
aud[21086]=16'h27d2;
aud[21087]=16'h27c1;
aud[21088]=16'h27b0;
aud[21089]=16'h279f;
aud[21090]=16'h278e;
aud[21091]=16'h277e;
aud[21092]=16'h276d;
aud[21093]=16'h275c;
aud[21094]=16'h274b;
aud[21095]=16'h273a;
aud[21096]=16'h2729;
aud[21097]=16'h2718;
aud[21098]=16'h2707;
aud[21099]=16'h26f6;
aud[21100]=16'h26e5;
aud[21101]=16'h26d4;
aud[21102]=16'h26c3;
aud[21103]=16'h26b2;
aud[21104]=16'h26a1;
aud[21105]=16'h2690;
aud[21106]=16'h267e;
aud[21107]=16'h266d;
aud[21108]=16'h265c;
aud[21109]=16'h264b;
aud[21110]=16'h263a;
aud[21111]=16'h2629;
aud[21112]=16'h2617;
aud[21113]=16'h2606;
aud[21114]=16'h25f5;
aud[21115]=16'h25e4;
aud[21116]=16'h25d2;
aud[21117]=16'h25c1;
aud[21118]=16'h25b0;
aud[21119]=16'h259e;
aud[21120]=16'h258d;
aud[21121]=16'h257c;
aud[21122]=16'h256a;
aud[21123]=16'h2559;
aud[21124]=16'h2547;
aud[21125]=16'h2536;
aud[21126]=16'h2524;
aud[21127]=16'h2513;
aud[21128]=16'h2501;
aud[21129]=16'h24f0;
aud[21130]=16'h24de;
aud[21131]=16'h24cd;
aud[21132]=16'h24bb;
aud[21133]=16'h24aa;
aud[21134]=16'h2498;
aud[21135]=16'h2487;
aud[21136]=16'h2475;
aud[21137]=16'h2463;
aud[21138]=16'h2452;
aud[21139]=16'h2440;
aud[21140]=16'h242e;
aud[21141]=16'h241d;
aud[21142]=16'h240b;
aud[21143]=16'h23f9;
aud[21144]=16'h23e7;
aud[21145]=16'h23d6;
aud[21146]=16'h23c4;
aud[21147]=16'h23b2;
aud[21148]=16'h23a0;
aud[21149]=16'h238e;
aud[21150]=16'h237d;
aud[21151]=16'h236b;
aud[21152]=16'h2359;
aud[21153]=16'h2347;
aud[21154]=16'h2335;
aud[21155]=16'h2323;
aud[21156]=16'h2311;
aud[21157]=16'h22ff;
aud[21158]=16'h22ed;
aud[21159]=16'h22db;
aud[21160]=16'h22c9;
aud[21161]=16'h22b7;
aud[21162]=16'h22a5;
aud[21163]=16'h2293;
aud[21164]=16'h2281;
aud[21165]=16'h226f;
aud[21166]=16'h225d;
aud[21167]=16'h224b;
aud[21168]=16'h2239;
aud[21169]=16'h2227;
aud[21170]=16'h2215;
aud[21171]=16'h2202;
aud[21172]=16'h21f0;
aud[21173]=16'h21de;
aud[21174]=16'h21cc;
aud[21175]=16'h21ba;
aud[21176]=16'h21a7;
aud[21177]=16'h2195;
aud[21178]=16'h2183;
aud[21179]=16'h2171;
aud[21180]=16'h215e;
aud[21181]=16'h214c;
aud[21182]=16'h213a;
aud[21183]=16'h2127;
aud[21184]=16'h2115;
aud[21185]=16'h2103;
aud[21186]=16'h20f0;
aud[21187]=16'h20de;
aud[21188]=16'h20cb;
aud[21189]=16'h20b9;
aud[21190]=16'h20a7;
aud[21191]=16'h2094;
aud[21192]=16'h2082;
aud[21193]=16'h206f;
aud[21194]=16'h205d;
aud[21195]=16'h204a;
aud[21196]=16'h2038;
aud[21197]=16'h2025;
aud[21198]=16'h2013;
aud[21199]=16'h2000;
aud[21200]=16'h1fed;
aud[21201]=16'h1fdb;
aud[21202]=16'h1fc8;
aud[21203]=16'h1fb6;
aud[21204]=16'h1fa3;
aud[21205]=16'h1f90;
aud[21206]=16'h1f7e;
aud[21207]=16'h1f6b;
aud[21208]=16'h1f58;
aud[21209]=16'h1f46;
aud[21210]=16'h1f33;
aud[21211]=16'h1f20;
aud[21212]=16'h1f0d;
aud[21213]=16'h1efb;
aud[21214]=16'h1ee8;
aud[21215]=16'h1ed5;
aud[21216]=16'h1ec2;
aud[21217]=16'h1eaf;
aud[21218]=16'h1e9d;
aud[21219]=16'h1e8a;
aud[21220]=16'h1e77;
aud[21221]=16'h1e64;
aud[21222]=16'h1e51;
aud[21223]=16'h1e3e;
aud[21224]=16'h1e2b;
aud[21225]=16'h1e18;
aud[21226]=16'h1e06;
aud[21227]=16'h1df3;
aud[21228]=16'h1de0;
aud[21229]=16'h1dcd;
aud[21230]=16'h1dba;
aud[21231]=16'h1da7;
aud[21232]=16'h1d94;
aud[21233]=16'h1d81;
aud[21234]=16'h1d6e;
aud[21235]=16'h1d5b;
aud[21236]=16'h1d47;
aud[21237]=16'h1d34;
aud[21238]=16'h1d21;
aud[21239]=16'h1d0e;
aud[21240]=16'h1cfb;
aud[21241]=16'h1ce8;
aud[21242]=16'h1cd5;
aud[21243]=16'h1cc2;
aud[21244]=16'h1cae;
aud[21245]=16'h1c9b;
aud[21246]=16'h1c88;
aud[21247]=16'h1c75;
aud[21248]=16'h1c62;
aud[21249]=16'h1c4e;
aud[21250]=16'h1c3b;
aud[21251]=16'h1c28;
aud[21252]=16'h1c15;
aud[21253]=16'h1c01;
aud[21254]=16'h1bee;
aud[21255]=16'h1bdb;
aud[21256]=16'h1bc8;
aud[21257]=16'h1bb4;
aud[21258]=16'h1ba1;
aud[21259]=16'h1b8d;
aud[21260]=16'h1b7a;
aud[21261]=16'h1b67;
aud[21262]=16'h1b53;
aud[21263]=16'h1b40;
aud[21264]=16'h1b2d;
aud[21265]=16'h1b19;
aud[21266]=16'h1b06;
aud[21267]=16'h1af2;
aud[21268]=16'h1adf;
aud[21269]=16'h1acb;
aud[21270]=16'h1ab8;
aud[21271]=16'h1aa4;
aud[21272]=16'h1a91;
aud[21273]=16'h1a7d;
aud[21274]=16'h1a6a;
aud[21275]=16'h1a56;
aud[21276]=16'h1a43;
aud[21277]=16'h1a2f;
aud[21278]=16'h1a1c;
aud[21279]=16'h1a08;
aud[21280]=16'h19f4;
aud[21281]=16'h19e1;
aud[21282]=16'h19cd;
aud[21283]=16'h19ba;
aud[21284]=16'h19a6;
aud[21285]=16'h1992;
aud[21286]=16'h197f;
aud[21287]=16'h196b;
aud[21288]=16'h1957;
aud[21289]=16'h1943;
aud[21290]=16'h1930;
aud[21291]=16'h191c;
aud[21292]=16'h1908;
aud[21293]=16'h18f5;
aud[21294]=16'h18e1;
aud[21295]=16'h18cd;
aud[21296]=16'h18b9;
aud[21297]=16'h18a5;
aud[21298]=16'h1892;
aud[21299]=16'h187e;
aud[21300]=16'h186a;
aud[21301]=16'h1856;
aud[21302]=16'h1842;
aud[21303]=16'h182f;
aud[21304]=16'h181b;
aud[21305]=16'h1807;
aud[21306]=16'h17f3;
aud[21307]=16'h17df;
aud[21308]=16'h17cb;
aud[21309]=16'h17b7;
aud[21310]=16'h17a3;
aud[21311]=16'h178f;
aud[21312]=16'h177b;
aud[21313]=16'h1767;
aud[21314]=16'h1753;
aud[21315]=16'h1740;
aud[21316]=16'h172c;
aud[21317]=16'h1718;
aud[21318]=16'h1704;
aud[21319]=16'h16f0;
aud[21320]=16'h16db;
aud[21321]=16'h16c7;
aud[21322]=16'h16b3;
aud[21323]=16'h169f;
aud[21324]=16'h168b;
aud[21325]=16'h1677;
aud[21326]=16'h1663;
aud[21327]=16'h164f;
aud[21328]=16'h163b;
aud[21329]=16'h1627;
aud[21330]=16'h1613;
aud[21331]=16'h15ff;
aud[21332]=16'h15ea;
aud[21333]=16'h15d6;
aud[21334]=16'h15c2;
aud[21335]=16'h15ae;
aud[21336]=16'h159a;
aud[21337]=16'h1586;
aud[21338]=16'h1571;
aud[21339]=16'h155d;
aud[21340]=16'h1549;
aud[21341]=16'h1535;
aud[21342]=16'h1520;
aud[21343]=16'h150c;
aud[21344]=16'h14f8;
aud[21345]=16'h14e4;
aud[21346]=16'h14cf;
aud[21347]=16'h14bb;
aud[21348]=16'h14a7;
aud[21349]=16'h1492;
aud[21350]=16'h147e;
aud[21351]=16'h146a;
aud[21352]=16'h1455;
aud[21353]=16'h1441;
aud[21354]=16'h142d;
aud[21355]=16'h1418;
aud[21356]=16'h1404;
aud[21357]=16'h13f0;
aud[21358]=16'h13db;
aud[21359]=16'h13c7;
aud[21360]=16'h13b3;
aud[21361]=16'h139e;
aud[21362]=16'h138a;
aud[21363]=16'h1375;
aud[21364]=16'h1361;
aud[21365]=16'h134c;
aud[21366]=16'h1338;
aud[21367]=16'h1323;
aud[21368]=16'h130f;
aud[21369]=16'h12fb;
aud[21370]=16'h12e6;
aud[21371]=16'h12d2;
aud[21372]=16'h12bd;
aud[21373]=16'h12a9;
aud[21374]=16'h1294;
aud[21375]=16'h127f;
aud[21376]=16'h126b;
aud[21377]=16'h1256;
aud[21378]=16'h1242;
aud[21379]=16'h122d;
aud[21380]=16'h1219;
aud[21381]=16'h1204;
aud[21382]=16'h11f0;
aud[21383]=16'h11db;
aud[21384]=16'h11c6;
aud[21385]=16'h11b2;
aud[21386]=16'h119d;
aud[21387]=16'h1189;
aud[21388]=16'h1174;
aud[21389]=16'h115f;
aud[21390]=16'h114b;
aud[21391]=16'h1136;
aud[21392]=16'h1121;
aud[21393]=16'h110d;
aud[21394]=16'h10f8;
aud[21395]=16'h10e3;
aud[21396]=16'h10cf;
aud[21397]=16'h10ba;
aud[21398]=16'h10a5;
aud[21399]=16'h1090;
aud[21400]=16'h107c;
aud[21401]=16'h1067;
aud[21402]=16'h1052;
aud[21403]=16'h103e;
aud[21404]=16'h1029;
aud[21405]=16'h1014;
aud[21406]=16'hfff;
aud[21407]=16'hfeb;
aud[21408]=16'hfd6;
aud[21409]=16'hfc1;
aud[21410]=16'hfac;
aud[21411]=16'hf97;
aud[21412]=16'hf83;
aud[21413]=16'hf6e;
aud[21414]=16'hf59;
aud[21415]=16'hf44;
aud[21416]=16'hf2f;
aud[21417]=16'hf1a;
aud[21418]=16'hf06;
aud[21419]=16'hef1;
aud[21420]=16'hedc;
aud[21421]=16'hec7;
aud[21422]=16'heb2;
aud[21423]=16'he9d;
aud[21424]=16'he88;
aud[21425]=16'he74;
aud[21426]=16'he5f;
aud[21427]=16'he4a;
aud[21428]=16'he35;
aud[21429]=16'he20;
aud[21430]=16'he0b;
aud[21431]=16'hdf6;
aud[21432]=16'hde1;
aud[21433]=16'hdcc;
aud[21434]=16'hdb7;
aud[21435]=16'hda2;
aud[21436]=16'hd8d;
aud[21437]=16'hd78;
aud[21438]=16'hd63;
aud[21439]=16'hd4e;
aud[21440]=16'hd39;
aud[21441]=16'hd24;
aud[21442]=16'hd0f;
aud[21443]=16'hcfa;
aud[21444]=16'hce5;
aud[21445]=16'hcd0;
aud[21446]=16'hcbb;
aud[21447]=16'hca6;
aud[21448]=16'hc91;
aud[21449]=16'hc7c;
aud[21450]=16'hc67;
aud[21451]=16'hc52;
aud[21452]=16'hc3d;
aud[21453]=16'hc28;
aud[21454]=16'hc13;
aud[21455]=16'hbfe;
aud[21456]=16'hbe9;
aud[21457]=16'hbd4;
aud[21458]=16'hbbf;
aud[21459]=16'hbaa;
aud[21460]=16'hb95;
aud[21461]=16'hb80;
aud[21462]=16'hb6a;
aud[21463]=16'hb55;
aud[21464]=16'hb40;
aud[21465]=16'hb2b;
aud[21466]=16'hb16;
aud[21467]=16'hb01;
aud[21468]=16'haec;
aud[21469]=16'had7;
aud[21470]=16'hac1;
aud[21471]=16'haac;
aud[21472]=16'ha97;
aud[21473]=16'ha82;
aud[21474]=16'ha6d;
aud[21475]=16'ha58;
aud[21476]=16'ha43;
aud[21477]=16'ha2d;
aud[21478]=16'ha18;
aud[21479]=16'ha03;
aud[21480]=16'h9ee;
aud[21481]=16'h9d9;
aud[21482]=16'h9c3;
aud[21483]=16'h9ae;
aud[21484]=16'h999;
aud[21485]=16'h984;
aud[21486]=16'h96f;
aud[21487]=16'h959;
aud[21488]=16'h944;
aud[21489]=16'h92f;
aud[21490]=16'h91a;
aud[21491]=16'h905;
aud[21492]=16'h8ef;
aud[21493]=16'h8da;
aud[21494]=16'h8c5;
aud[21495]=16'h8b0;
aud[21496]=16'h89a;
aud[21497]=16'h885;
aud[21498]=16'h870;
aud[21499]=16'h85b;
aud[21500]=16'h845;
aud[21501]=16'h830;
aud[21502]=16'h81b;
aud[21503]=16'h805;
aud[21504]=16'h7f0;
aud[21505]=16'h7db;
aud[21506]=16'h7c6;
aud[21507]=16'h7b0;
aud[21508]=16'h79b;
aud[21509]=16'h786;
aud[21510]=16'h770;
aud[21511]=16'h75b;
aud[21512]=16'h746;
aud[21513]=16'h731;
aud[21514]=16'h71b;
aud[21515]=16'h706;
aud[21516]=16'h6f1;
aud[21517]=16'h6db;
aud[21518]=16'h6c6;
aud[21519]=16'h6b1;
aud[21520]=16'h69b;
aud[21521]=16'h686;
aud[21522]=16'h671;
aud[21523]=16'h65b;
aud[21524]=16'h646;
aud[21525]=16'h631;
aud[21526]=16'h61b;
aud[21527]=16'h606;
aud[21528]=16'h5f1;
aud[21529]=16'h5db;
aud[21530]=16'h5c6;
aud[21531]=16'h5b0;
aud[21532]=16'h59b;
aud[21533]=16'h586;
aud[21534]=16'h570;
aud[21535]=16'h55b;
aud[21536]=16'h546;
aud[21537]=16'h530;
aud[21538]=16'h51b;
aud[21539]=16'h505;
aud[21540]=16'h4f0;
aud[21541]=16'h4db;
aud[21542]=16'h4c5;
aud[21543]=16'h4b0;
aud[21544]=16'h49b;
aud[21545]=16'h485;
aud[21546]=16'h470;
aud[21547]=16'h45a;
aud[21548]=16'h445;
aud[21549]=16'h430;
aud[21550]=16'h41a;
aud[21551]=16'h405;
aud[21552]=16'h3ef;
aud[21553]=16'h3da;
aud[21554]=16'h3c5;
aud[21555]=16'h3af;
aud[21556]=16'h39a;
aud[21557]=16'h384;
aud[21558]=16'h36f;
aud[21559]=16'h359;
aud[21560]=16'h344;
aud[21561]=16'h32f;
aud[21562]=16'h319;
aud[21563]=16'h304;
aud[21564]=16'h2ee;
aud[21565]=16'h2d9;
aud[21566]=16'h2c4;
aud[21567]=16'h2ae;
aud[21568]=16'h299;
aud[21569]=16'h283;
aud[21570]=16'h26e;
aud[21571]=16'h258;
aud[21572]=16'h243;
aud[21573]=16'h22e;
aud[21574]=16'h218;
aud[21575]=16'h203;
aud[21576]=16'h1ed;
aud[21577]=16'h1d8;
aud[21578]=16'h1c2;
aud[21579]=16'h1ad;
aud[21580]=16'h197;
aud[21581]=16'h182;
aud[21582]=16'h16d;
aud[21583]=16'h157;
aud[21584]=16'h142;
aud[21585]=16'h12c;
aud[21586]=16'h117;
aud[21587]=16'h101;
aud[21588]=16'hec;
aud[21589]=16'hd6;
aud[21590]=16'hc1;
aud[21591]=16'hac;
aud[21592]=16'h96;
aud[21593]=16'h81;
aud[21594]=16'h6b;
aud[21595]=16'h56;
aud[21596]=16'h40;
aud[21597]=16'h2b;
aud[21598]=16'h15;
aud[21599]=16'h0;
aud[21600]=16'hffeb;
aud[21601]=16'hffd5;
aud[21602]=16'hffc0;
aud[21603]=16'hffaa;
aud[21604]=16'hff95;
aud[21605]=16'hff7f;
aud[21606]=16'hff6a;
aud[21607]=16'hff54;
aud[21608]=16'hff3f;
aud[21609]=16'hff2a;
aud[21610]=16'hff14;
aud[21611]=16'hfeff;
aud[21612]=16'hfee9;
aud[21613]=16'hfed4;
aud[21614]=16'hfebe;
aud[21615]=16'hfea9;
aud[21616]=16'hfe93;
aud[21617]=16'hfe7e;
aud[21618]=16'hfe69;
aud[21619]=16'hfe53;
aud[21620]=16'hfe3e;
aud[21621]=16'hfe28;
aud[21622]=16'hfe13;
aud[21623]=16'hfdfd;
aud[21624]=16'hfde8;
aud[21625]=16'hfdd2;
aud[21626]=16'hfdbd;
aud[21627]=16'hfda8;
aud[21628]=16'hfd92;
aud[21629]=16'hfd7d;
aud[21630]=16'hfd67;
aud[21631]=16'hfd52;
aud[21632]=16'hfd3c;
aud[21633]=16'hfd27;
aud[21634]=16'hfd12;
aud[21635]=16'hfcfc;
aud[21636]=16'hfce7;
aud[21637]=16'hfcd1;
aud[21638]=16'hfcbc;
aud[21639]=16'hfca7;
aud[21640]=16'hfc91;
aud[21641]=16'hfc7c;
aud[21642]=16'hfc66;
aud[21643]=16'hfc51;
aud[21644]=16'hfc3b;
aud[21645]=16'hfc26;
aud[21646]=16'hfc11;
aud[21647]=16'hfbfb;
aud[21648]=16'hfbe6;
aud[21649]=16'hfbd0;
aud[21650]=16'hfbbb;
aud[21651]=16'hfba6;
aud[21652]=16'hfb90;
aud[21653]=16'hfb7b;
aud[21654]=16'hfb65;
aud[21655]=16'hfb50;
aud[21656]=16'hfb3b;
aud[21657]=16'hfb25;
aud[21658]=16'hfb10;
aud[21659]=16'hfafb;
aud[21660]=16'hfae5;
aud[21661]=16'hfad0;
aud[21662]=16'hfaba;
aud[21663]=16'hfaa5;
aud[21664]=16'hfa90;
aud[21665]=16'hfa7a;
aud[21666]=16'hfa65;
aud[21667]=16'hfa50;
aud[21668]=16'hfa3a;
aud[21669]=16'hfa25;
aud[21670]=16'hfa0f;
aud[21671]=16'hf9fa;
aud[21672]=16'hf9e5;
aud[21673]=16'hf9cf;
aud[21674]=16'hf9ba;
aud[21675]=16'hf9a5;
aud[21676]=16'hf98f;
aud[21677]=16'hf97a;
aud[21678]=16'hf965;
aud[21679]=16'hf94f;
aud[21680]=16'hf93a;
aud[21681]=16'hf925;
aud[21682]=16'hf90f;
aud[21683]=16'hf8fa;
aud[21684]=16'hf8e5;
aud[21685]=16'hf8cf;
aud[21686]=16'hf8ba;
aud[21687]=16'hf8a5;
aud[21688]=16'hf890;
aud[21689]=16'hf87a;
aud[21690]=16'hf865;
aud[21691]=16'hf850;
aud[21692]=16'hf83a;
aud[21693]=16'hf825;
aud[21694]=16'hf810;
aud[21695]=16'hf7fb;
aud[21696]=16'hf7e5;
aud[21697]=16'hf7d0;
aud[21698]=16'hf7bb;
aud[21699]=16'hf7a5;
aud[21700]=16'hf790;
aud[21701]=16'hf77b;
aud[21702]=16'hf766;
aud[21703]=16'hf750;
aud[21704]=16'hf73b;
aud[21705]=16'hf726;
aud[21706]=16'hf711;
aud[21707]=16'hf6fb;
aud[21708]=16'hf6e6;
aud[21709]=16'hf6d1;
aud[21710]=16'hf6bc;
aud[21711]=16'hf6a7;
aud[21712]=16'hf691;
aud[21713]=16'hf67c;
aud[21714]=16'hf667;
aud[21715]=16'hf652;
aud[21716]=16'hf63d;
aud[21717]=16'hf627;
aud[21718]=16'hf612;
aud[21719]=16'hf5fd;
aud[21720]=16'hf5e8;
aud[21721]=16'hf5d3;
aud[21722]=16'hf5bd;
aud[21723]=16'hf5a8;
aud[21724]=16'hf593;
aud[21725]=16'hf57e;
aud[21726]=16'hf569;
aud[21727]=16'hf554;
aud[21728]=16'hf53f;
aud[21729]=16'hf529;
aud[21730]=16'hf514;
aud[21731]=16'hf4ff;
aud[21732]=16'hf4ea;
aud[21733]=16'hf4d5;
aud[21734]=16'hf4c0;
aud[21735]=16'hf4ab;
aud[21736]=16'hf496;
aud[21737]=16'hf480;
aud[21738]=16'hf46b;
aud[21739]=16'hf456;
aud[21740]=16'hf441;
aud[21741]=16'hf42c;
aud[21742]=16'hf417;
aud[21743]=16'hf402;
aud[21744]=16'hf3ed;
aud[21745]=16'hf3d8;
aud[21746]=16'hf3c3;
aud[21747]=16'hf3ae;
aud[21748]=16'hf399;
aud[21749]=16'hf384;
aud[21750]=16'hf36f;
aud[21751]=16'hf35a;
aud[21752]=16'hf345;
aud[21753]=16'hf330;
aud[21754]=16'hf31b;
aud[21755]=16'hf306;
aud[21756]=16'hf2f1;
aud[21757]=16'hf2dc;
aud[21758]=16'hf2c7;
aud[21759]=16'hf2b2;
aud[21760]=16'hf29d;
aud[21761]=16'hf288;
aud[21762]=16'hf273;
aud[21763]=16'hf25e;
aud[21764]=16'hf249;
aud[21765]=16'hf234;
aud[21766]=16'hf21f;
aud[21767]=16'hf20a;
aud[21768]=16'hf1f5;
aud[21769]=16'hf1e0;
aud[21770]=16'hf1cb;
aud[21771]=16'hf1b6;
aud[21772]=16'hf1a1;
aud[21773]=16'hf18c;
aud[21774]=16'hf178;
aud[21775]=16'hf163;
aud[21776]=16'hf14e;
aud[21777]=16'hf139;
aud[21778]=16'hf124;
aud[21779]=16'hf10f;
aud[21780]=16'hf0fa;
aud[21781]=16'hf0e6;
aud[21782]=16'hf0d1;
aud[21783]=16'hf0bc;
aud[21784]=16'hf0a7;
aud[21785]=16'hf092;
aud[21786]=16'hf07d;
aud[21787]=16'hf069;
aud[21788]=16'hf054;
aud[21789]=16'hf03f;
aud[21790]=16'hf02a;
aud[21791]=16'hf015;
aud[21792]=16'hf001;
aud[21793]=16'hefec;
aud[21794]=16'hefd7;
aud[21795]=16'hefc2;
aud[21796]=16'hefae;
aud[21797]=16'hef99;
aud[21798]=16'hef84;
aud[21799]=16'hef70;
aud[21800]=16'hef5b;
aud[21801]=16'hef46;
aud[21802]=16'hef31;
aud[21803]=16'hef1d;
aud[21804]=16'hef08;
aud[21805]=16'heef3;
aud[21806]=16'heedf;
aud[21807]=16'heeca;
aud[21808]=16'heeb5;
aud[21809]=16'heea1;
aud[21810]=16'hee8c;
aud[21811]=16'hee77;
aud[21812]=16'hee63;
aud[21813]=16'hee4e;
aud[21814]=16'hee3a;
aud[21815]=16'hee25;
aud[21816]=16'hee10;
aud[21817]=16'hedfc;
aud[21818]=16'hede7;
aud[21819]=16'hedd3;
aud[21820]=16'hedbe;
aud[21821]=16'hedaa;
aud[21822]=16'hed95;
aud[21823]=16'hed81;
aud[21824]=16'hed6c;
aud[21825]=16'hed57;
aud[21826]=16'hed43;
aud[21827]=16'hed2e;
aud[21828]=16'hed1a;
aud[21829]=16'hed05;
aud[21830]=16'hecf1;
aud[21831]=16'hecdd;
aud[21832]=16'hecc8;
aud[21833]=16'hecb4;
aud[21834]=16'hec9f;
aud[21835]=16'hec8b;
aud[21836]=16'hec76;
aud[21837]=16'hec62;
aud[21838]=16'hec4d;
aud[21839]=16'hec39;
aud[21840]=16'hec25;
aud[21841]=16'hec10;
aud[21842]=16'hebfc;
aud[21843]=16'hebe8;
aud[21844]=16'hebd3;
aud[21845]=16'hebbf;
aud[21846]=16'hebab;
aud[21847]=16'heb96;
aud[21848]=16'heb82;
aud[21849]=16'heb6e;
aud[21850]=16'heb59;
aud[21851]=16'heb45;
aud[21852]=16'heb31;
aud[21853]=16'heb1c;
aud[21854]=16'heb08;
aud[21855]=16'heaf4;
aud[21856]=16'heae0;
aud[21857]=16'heacb;
aud[21858]=16'heab7;
aud[21859]=16'heaa3;
aud[21860]=16'hea8f;
aud[21861]=16'hea7a;
aud[21862]=16'hea66;
aud[21863]=16'hea52;
aud[21864]=16'hea3e;
aud[21865]=16'hea2a;
aud[21866]=16'hea16;
aud[21867]=16'hea01;
aud[21868]=16'he9ed;
aud[21869]=16'he9d9;
aud[21870]=16'he9c5;
aud[21871]=16'he9b1;
aud[21872]=16'he99d;
aud[21873]=16'he989;
aud[21874]=16'he975;
aud[21875]=16'he961;
aud[21876]=16'he94d;
aud[21877]=16'he939;
aud[21878]=16'he925;
aud[21879]=16'he910;
aud[21880]=16'he8fc;
aud[21881]=16'he8e8;
aud[21882]=16'he8d4;
aud[21883]=16'he8c0;
aud[21884]=16'he8ad;
aud[21885]=16'he899;
aud[21886]=16'he885;
aud[21887]=16'he871;
aud[21888]=16'he85d;
aud[21889]=16'he849;
aud[21890]=16'he835;
aud[21891]=16'he821;
aud[21892]=16'he80d;
aud[21893]=16'he7f9;
aud[21894]=16'he7e5;
aud[21895]=16'he7d1;
aud[21896]=16'he7be;
aud[21897]=16'he7aa;
aud[21898]=16'he796;
aud[21899]=16'he782;
aud[21900]=16'he76e;
aud[21901]=16'he75b;
aud[21902]=16'he747;
aud[21903]=16'he733;
aud[21904]=16'he71f;
aud[21905]=16'he70b;
aud[21906]=16'he6f8;
aud[21907]=16'he6e4;
aud[21908]=16'he6d0;
aud[21909]=16'he6bd;
aud[21910]=16'he6a9;
aud[21911]=16'he695;
aud[21912]=16'he681;
aud[21913]=16'he66e;
aud[21914]=16'he65a;
aud[21915]=16'he646;
aud[21916]=16'he633;
aud[21917]=16'he61f;
aud[21918]=16'he60c;
aud[21919]=16'he5f8;
aud[21920]=16'he5e4;
aud[21921]=16'he5d1;
aud[21922]=16'he5bd;
aud[21923]=16'he5aa;
aud[21924]=16'he596;
aud[21925]=16'he583;
aud[21926]=16'he56f;
aud[21927]=16'he55c;
aud[21928]=16'he548;
aud[21929]=16'he535;
aud[21930]=16'he521;
aud[21931]=16'he50e;
aud[21932]=16'he4fa;
aud[21933]=16'he4e7;
aud[21934]=16'he4d3;
aud[21935]=16'he4c0;
aud[21936]=16'he4ad;
aud[21937]=16'he499;
aud[21938]=16'he486;
aud[21939]=16'he473;
aud[21940]=16'he45f;
aud[21941]=16'he44c;
aud[21942]=16'he438;
aud[21943]=16'he425;
aud[21944]=16'he412;
aud[21945]=16'he3ff;
aud[21946]=16'he3eb;
aud[21947]=16'he3d8;
aud[21948]=16'he3c5;
aud[21949]=16'he3b2;
aud[21950]=16'he39e;
aud[21951]=16'he38b;
aud[21952]=16'he378;
aud[21953]=16'he365;
aud[21954]=16'he352;
aud[21955]=16'he33e;
aud[21956]=16'he32b;
aud[21957]=16'he318;
aud[21958]=16'he305;
aud[21959]=16'he2f2;
aud[21960]=16'he2df;
aud[21961]=16'he2cc;
aud[21962]=16'he2b9;
aud[21963]=16'he2a5;
aud[21964]=16'he292;
aud[21965]=16'he27f;
aud[21966]=16'he26c;
aud[21967]=16'he259;
aud[21968]=16'he246;
aud[21969]=16'he233;
aud[21970]=16'he220;
aud[21971]=16'he20d;
aud[21972]=16'he1fa;
aud[21973]=16'he1e8;
aud[21974]=16'he1d5;
aud[21975]=16'he1c2;
aud[21976]=16'he1af;
aud[21977]=16'he19c;
aud[21978]=16'he189;
aud[21979]=16'he176;
aud[21980]=16'he163;
aud[21981]=16'he151;
aud[21982]=16'he13e;
aud[21983]=16'he12b;
aud[21984]=16'he118;
aud[21985]=16'he105;
aud[21986]=16'he0f3;
aud[21987]=16'he0e0;
aud[21988]=16'he0cd;
aud[21989]=16'he0ba;
aud[21990]=16'he0a8;
aud[21991]=16'he095;
aud[21992]=16'he082;
aud[21993]=16'he070;
aud[21994]=16'he05d;
aud[21995]=16'he04a;
aud[21996]=16'he038;
aud[21997]=16'he025;
aud[21998]=16'he013;
aud[21999]=16'he000;
aud[22000]=16'hdfed;
aud[22001]=16'hdfdb;
aud[22002]=16'hdfc8;
aud[22003]=16'hdfb6;
aud[22004]=16'hdfa3;
aud[22005]=16'hdf91;
aud[22006]=16'hdf7e;
aud[22007]=16'hdf6c;
aud[22008]=16'hdf59;
aud[22009]=16'hdf47;
aud[22010]=16'hdf35;
aud[22011]=16'hdf22;
aud[22012]=16'hdf10;
aud[22013]=16'hdefd;
aud[22014]=16'hdeeb;
aud[22015]=16'hded9;
aud[22016]=16'hdec6;
aud[22017]=16'hdeb4;
aud[22018]=16'hdea2;
aud[22019]=16'hde8f;
aud[22020]=16'hde7d;
aud[22021]=16'hde6b;
aud[22022]=16'hde59;
aud[22023]=16'hde46;
aud[22024]=16'hde34;
aud[22025]=16'hde22;
aud[22026]=16'hde10;
aud[22027]=16'hddfe;
aud[22028]=16'hddeb;
aud[22029]=16'hddd9;
aud[22030]=16'hddc7;
aud[22031]=16'hddb5;
aud[22032]=16'hdda3;
aud[22033]=16'hdd91;
aud[22034]=16'hdd7f;
aud[22035]=16'hdd6d;
aud[22036]=16'hdd5b;
aud[22037]=16'hdd49;
aud[22038]=16'hdd37;
aud[22039]=16'hdd25;
aud[22040]=16'hdd13;
aud[22041]=16'hdd01;
aud[22042]=16'hdcef;
aud[22043]=16'hdcdd;
aud[22044]=16'hdccb;
aud[22045]=16'hdcb9;
aud[22046]=16'hdca7;
aud[22047]=16'hdc95;
aud[22048]=16'hdc83;
aud[22049]=16'hdc72;
aud[22050]=16'hdc60;
aud[22051]=16'hdc4e;
aud[22052]=16'hdc3c;
aud[22053]=16'hdc2a;
aud[22054]=16'hdc19;
aud[22055]=16'hdc07;
aud[22056]=16'hdbf5;
aud[22057]=16'hdbe3;
aud[22058]=16'hdbd2;
aud[22059]=16'hdbc0;
aud[22060]=16'hdbae;
aud[22061]=16'hdb9d;
aud[22062]=16'hdb8b;
aud[22063]=16'hdb79;
aud[22064]=16'hdb68;
aud[22065]=16'hdb56;
aud[22066]=16'hdb45;
aud[22067]=16'hdb33;
aud[22068]=16'hdb22;
aud[22069]=16'hdb10;
aud[22070]=16'hdaff;
aud[22071]=16'hdaed;
aud[22072]=16'hdadc;
aud[22073]=16'hdaca;
aud[22074]=16'hdab9;
aud[22075]=16'hdaa7;
aud[22076]=16'hda96;
aud[22077]=16'hda84;
aud[22078]=16'hda73;
aud[22079]=16'hda62;
aud[22080]=16'hda50;
aud[22081]=16'hda3f;
aud[22082]=16'hda2e;
aud[22083]=16'hda1c;
aud[22084]=16'hda0b;
aud[22085]=16'hd9fa;
aud[22086]=16'hd9e9;
aud[22087]=16'hd9d7;
aud[22088]=16'hd9c6;
aud[22089]=16'hd9b5;
aud[22090]=16'hd9a4;
aud[22091]=16'hd993;
aud[22092]=16'hd982;
aud[22093]=16'hd970;
aud[22094]=16'hd95f;
aud[22095]=16'hd94e;
aud[22096]=16'hd93d;
aud[22097]=16'hd92c;
aud[22098]=16'hd91b;
aud[22099]=16'hd90a;
aud[22100]=16'hd8f9;
aud[22101]=16'hd8e8;
aud[22102]=16'hd8d7;
aud[22103]=16'hd8c6;
aud[22104]=16'hd8b5;
aud[22105]=16'hd8a4;
aud[22106]=16'hd893;
aud[22107]=16'hd882;
aud[22108]=16'hd872;
aud[22109]=16'hd861;
aud[22110]=16'hd850;
aud[22111]=16'hd83f;
aud[22112]=16'hd82e;
aud[22113]=16'hd81e;
aud[22114]=16'hd80d;
aud[22115]=16'hd7fc;
aud[22116]=16'hd7eb;
aud[22117]=16'hd7db;
aud[22118]=16'hd7ca;
aud[22119]=16'hd7b9;
aud[22120]=16'hd7a9;
aud[22121]=16'hd798;
aud[22122]=16'hd787;
aud[22123]=16'hd777;
aud[22124]=16'hd766;
aud[22125]=16'hd756;
aud[22126]=16'hd745;
aud[22127]=16'hd734;
aud[22128]=16'hd724;
aud[22129]=16'hd713;
aud[22130]=16'hd703;
aud[22131]=16'hd6f2;
aud[22132]=16'hd6e2;
aud[22133]=16'hd6d2;
aud[22134]=16'hd6c1;
aud[22135]=16'hd6b1;
aud[22136]=16'hd6a0;
aud[22137]=16'hd690;
aud[22138]=16'hd680;
aud[22139]=16'hd66f;
aud[22140]=16'hd65f;
aud[22141]=16'hd64f;
aud[22142]=16'hd63f;
aud[22143]=16'hd62e;
aud[22144]=16'hd61e;
aud[22145]=16'hd60e;
aud[22146]=16'hd5fe;
aud[22147]=16'hd5ee;
aud[22148]=16'hd5dd;
aud[22149]=16'hd5cd;
aud[22150]=16'hd5bd;
aud[22151]=16'hd5ad;
aud[22152]=16'hd59d;
aud[22153]=16'hd58d;
aud[22154]=16'hd57d;
aud[22155]=16'hd56d;
aud[22156]=16'hd55d;
aud[22157]=16'hd54d;
aud[22158]=16'hd53d;
aud[22159]=16'hd52d;
aud[22160]=16'hd51d;
aud[22161]=16'hd50d;
aud[22162]=16'hd4fd;
aud[22163]=16'hd4ed;
aud[22164]=16'hd4de;
aud[22165]=16'hd4ce;
aud[22166]=16'hd4be;
aud[22167]=16'hd4ae;
aud[22168]=16'hd49e;
aud[22169]=16'hd48f;
aud[22170]=16'hd47f;
aud[22171]=16'hd46f;
aud[22172]=16'hd45f;
aud[22173]=16'hd450;
aud[22174]=16'hd440;
aud[22175]=16'hd430;
aud[22176]=16'hd421;
aud[22177]=16'hd411;
aud[22178]=16'hd402;
aud[22179]=16'hd3f2;
aud[22180]=16'hd3e2;
aud[22181]=16'hd3d3;
aud[22182]=16'hd3c3;
aud[22183]=16'hd3b4;
aud[22184]=16'hd3a4;
aud[22185]=16'hd395;
aud[22186]=16'hd386;
aud[22187]=16'hd376;
aud[22188]=16'hd367;
aud[22189]=16'hd357;
aud[22190]=16'hd348;
aud[22191]=16'hd339;
aud[22192]=16'hd329;
aud[22193]=16'hd31a;
aud[22194]=16'hd30b;
aud[22195]=16'hd2fc;
aud[22196]=16'hd2ec;
aud[22197]=16'hd2dd;
aud[22198]=16'hd2ce;
aud[22199]=16'hd2bf;
aud[22200]=16'hd2b0;
aud[22201]=16'hd2a0;
aud[22202]=16'hd291;
aud[22203]=16'hd282;
aud[22204]=16'hd273;
aud[22205]=16'hd264;
aud[22206]=16'hd255;
aud[22207]=16'hd246;
aud[22208]=16'hd237;
aud[22209]=16'hd228;
aud[22210]=16'hd219;
aud[22211]=16'hd20a;
aud[22212]=16'hd1fb;
aud[22213]=16'hd1ec;
aud[22214]=16'hd1de;
aud[22215]=16'hd1cf;
aud[22216]=16'hd1c0;
aud[22217]=16'hd1b1;
aud[22218]=16'hd1a2;
aud[22219]=16'hd193;
aud[22220]=16'hd185;
aud[22221]=16'hd176;
aud[22222]=16'hd167;
aud[22223]=16'hd159;
aud[22224]=16'hd14a;
aud[22225]=16'hd13b;
aud[22226]=16'hd12d;
aud[22227]=16'hd11e;
aud[22228]=16'hd10f;
aud[22229]=16'hd101;
aud[22230]=16'hd0f2;
aud[22231]=16'hd0e4;
aud[22232]=16'hd0d5;
aud[22233]=16'hd0c7;
aud[22234]=16'hd0b8;
aud[22235]=16'hd0aa;
aud[22236]=16'hd09b;
aud[22237]=16'hd08d;
aud[22238]=16'hd07f;
aud[22239]=16'hd070;
aud[22240]=16'hd062;
aud[22241]=16'hd054;
aud[22242]=16'hd045;
aud[22243]=16'hd037;
aud[22244]=16'hd029;
aud[22245]=16'hd01b;
aud[22246]=16'hd00c;
aud[22247]=16'hcffe;
aud[22248]=16'hcff0;
aud[22249]=16'hcfe2;
aud[22250]=16'hcfd4;
aud[22251]=16'hcfc6;
aud[22252]=16'hcfb8;
aud[22253]=16'hcfa9;
aud[22254]=16'hcf9b;
aud[22255]=16'hcf8d;
aud[22256]=16'hcf7f;
aud[22257]=16'hcf71;
aud[22258]=16'hcf63;
aud[22259]=16'hcf56;
aud[22260]=16'hcf48;
aud[22261]=16'hcf3a;
aud[22262]=16'hcf2c;
aud[22263]=16'hcf1e;
aud[22264]=16'hcf10;
aud[22265]=16'hcf02;
aud[22266]=16'hcef5;
aud[22267]=16'hcee7;
aud[22268]=16'hced9;
aud[22269]=16'hcecb;
aud[22270]=16'hcebe;
aud[22271]=16'hceb0;
aud[22272]=16'hcea2;
aud[22273]=16'hce95;
aud[22274]=16'hce87;
aud[22275]=16'hce79;
aud[22276]=16'hce6c;
aud[22277]=16'hce5e;
aud[22278]=16'hce51;
aud[22279]=16'hce43;
aud[22280]=16'hce36;
aud[22281]=16'hce28;
aud[22282]=16'hce1b;
aud[22283]=16'hce0d;
aud[22284]=16'hce00;
aud[22285]=16'hcdf3;
aud[22286]=16'hcde5;
aud[22287]=16'hcdd8;
aud[22288]=16'hcdcb;
aud[22289]=16'hcdbd;
aud[22290]=16'hcdb0;
aud[22291]=16'hcda3;
aud[22292]=16'hcd96;
aud[22293]=16'hcd88;
aud[22294]=16'hcd7b;
aud[22295]=16'hcd6e;
aud[22296]=16'hcd61;
aud[22297]=16'hcd54;
aud[22298]=16'hcd47;
aud[22299]=16'hcd3a;
aud[22300]=16'hcd2d;
aud[22301]=16'hcd20;
aud[22302]=16'hcd13;
aud[22303]=16'hcd06;
aud[22304]=16'hccf9;
aud[22305]=16'hccec;
aud[22306]=16'hccdf;
aud[22307]=16'hccd2;
aud[22308]=16'hccc5;
aud[22309]=16'hccb8;
aud[22310]=16'hccab;
aud[22311]=16'hcc9f;
aud[22312]=16'hcc92;
aud[22313]=16'hcc85;
aud[22314]=16'hcc78;
aud[22315]=16'hcc6c;
aud[22316]=16'hcc5f;
aud[22317]=16'hcc52;
aud[22318]=16'hcc46;
aud[22319]=16'hcc39;
aud[22320]=16'hcc2c;
aud[22321]=16'hcc20;
aud[22322]=16'hcc13;
aud[22323]=16'hcc07;
aud[22324]=16'hcbfa;
aud[22325]=16'hcbee;
aud[22326]=16'hcbe1;
aud[22327]=16'hcbd5;
aud[22328]=16'hcbc9;
aud[22329]=16'hcbbc;
aud[22330]=16'hcbb0;
aud[22331]=16'hcba3;
aud[22332]=16'hcb97;
aud[22333]=16'hcb8b;
aud[22334]=16'hcb7f;
aud[22335]=16'hcb72;
aud[22336]=16'hcb66;
aud[22337]=16'hcb5a;
aud[22338]=16'hcb4e;
aud[22339]=16'hcb42;
aud[22340]=16'hcb35;
aud[22341]=16'hcb29;
aud[22342]=16'hcb1d;
aud[22343]=16'hcb11;
aud[22344]=16'hcb05;
aud[22345]=16'hcaf9;
aud[22346]=16'hcaed;
aud[22347]=16'hcae1;
aud[22348]=16'hcad5;
aud[22349]=16'hcac9;
aud[22350]=16'hcabd;
aud[22351]=16'hcab1;
aud[22352]=16'hcaa6;
aud[22353]=16'hca9a;
aud[22354]=16'hca8e;
aud[22355]=16'hca82;
aud[22356]=16'hca76;
aud[22357]=16'hca6b;
aud[22358]=16'hca5f;
aud[22359]=16'hca53;
aud[22360]=16'hca48;
aud[22361]=16'hca3c;
aud[22362]=16'hca30;
aud[22363]=16'hca25;
aud[22364]=16'hca19;
aud[22365]=16'hca0e;
aud[22366]=16'hca02;
aud[22367]=16'hc9f7;
aud[22368]=16'hc9eb;
aud[22369]=16'hc9e0;
aud[22370]=16'hc9d4;
aud[22371]=16'hc9c9;
aud[22372]=16'hc9bd;
aud[22373]=16'hc9b2;
aud[22374]=16'hc9a7;
aud[22375]=16'hc99b;
aud[22376]=16'hc990;
aud[22377]=16'hc985;
aud[22378]=16'hc97a;
aud[22379]=16'hc96e;
aud[22380]=16'hc963;
aud[22381]=16'hc958;
aud[22382]=16'hc94d;
aud[22383]=16'hc942;
aud[22384]=16'hc937;
aud[22385]=16'hc92c;
aud[22386]=16'hc920;
aud[22387]=16'hc915;
aud[22388]=16'hc90a;
aud[22389]=16'hc8ff;
aud[22390]=16'hc8f5;
aud[22391]=16'hc8ea;
aud[22392]=16'hc8df;
aud[22393]=16'hc8d4;
aud[22394]=16'hc8c9;
aud[22395]=16'hc8be;
aud[22396]=16'hc8b3;
aud[22397]=16'hc8a9;
aud[22398]=16'hc89e;
aud[22399]=16'hc893;
aud[22400]=16'hc888;
aud[22401]=16'hc87e;
aud[22402]=16'hc873;
aud[22403]=16'hc868;
aud[22404]=16'hc85e;
aud[22405]=16'hc853;
aud[22406]=16'hc849;
aud[22407]=16'hc83e;
aud[22408]=16'hc834;
aud[22409]=16'hc829;
aud[22410]=16'hc81f;
aud[22411]=16'hc814;
aud[22412]=16'hc80a;
aud[22413]=16'hc7ff;
aud[22414]=16'hc7f5;
aud[22415]=16'hc7eb;
aud[22416]=16'hc7e0;
aud[22417]=16'hc7d6;
aud[22418]=16'hc7cc;
aud[22419]=16'hc7c1;
aud[22420]=16'hc7b7;
aud[22421]=16'hc7ad;
aud[22422]=16'hc7a3;
aud[22423]=16'hc799;
aud[22424]=16'hc78f;
aud[22425]=16'hc785;
aud[22426]=16'hc77a;
aud[22427]=16'hc770;
aud[22428]=16'hc766;
aud[22429]=16'hc75c;
aud[22430]=16'hc752;
aud[22431]=16'hc748;
aud[22432]=16'hc73f;
aud[22433]=16'hc735;
aud[22434]=16'hc72b;
aud[22435]=16'hc721;
aud[22436]=16'hc717;
aud[22437]=16'hc70d;
aud[22438]=16'hc703;
aud[22439]=16'hc6fa;
aud[22440]=16'hc6f0;
aud[22441]=16'hc6e6;
aud[22442]=16'hc6dd;
aud[22443]=16'hc6d3;
aud[22444]=16'hc6c9;
aud[22445]=16'hc6c0;
aud[22446]=16'hc6b6;
aud[22447]=16'hc6ad;
aud[22448]=16'hc6a3;
aud[22449]=16'hc69a;
aud[22450]=16'hc690;
aud[22451]=16'hc687;
aud[22452]=16'hc67d;
aud[22453]=16'hc674;
aud[22454]=16'hc66b;
aud[22455]=16'hc661;
aud[22456]=16'hc658;
aud[22457]=16'hc64f;
aud[22458]=16'hc645;
aud[22459]=16'hc63c;
aud[22460]=16'hc633;
aud[22461]=16'hc62a;
aud[22462]=16'hc620;
aud[22463]=16'hc617;
aud[22464]=16'hc60e;
aud[22465]=16'hc605;
aud[22466]=16'hc5fc;
aud[22467]=16'hc5f3;
aud[22468]=16'hc5ea;
aud[22469]=16'hc5e1;
aud[22470]=16'hc5d8;
aud[22471]=16'hc5cf;
aud[22472]=16'hc5c6;
aud[22473]=16'hc5bd;
aud[22474]=16'hc5b4;
aud[22475]=16'hc5ac;
aud[22476]=16'hc5a3;
aud[22477]=16'hc59a;
aud[22478]=16'hc591;
aud[22479]=16'hc588;
aud[22480]=16'hc580;
aud[22481]=16'hc577;
aud[22482]=16'hc56e;
aud[22483]=16'hc566;
aud[22484]=16'hc55d;
aud[22485]=16'hc555;
aud[22486]=16'hc54c;
aud[22487]=16'hc544;
aud[22488]=16'hc53b;
aud[22489]=16'hc533;
aud[22490]=16'hc52a;
aud[22491]=16'hc522;
aud[22492]=16'hc519;
aud[22493]=16'hc511;
aud[22494]=16'hc509;
aud[22495]=16'hc500;
aud[22496]=16'hc4f8;
aud[22497]=16'hc4f0;
aud[22498]=16'hc4e7;
aud[22499]=16'hc4df;
aud[22500]=16'hc4d7;
aud[22501]=16'hc4cf;
aud[22502]=16'hc4c7;
aud[22503]=16'hc4bf;
aud[22504]=16'hc4b6;
aud[22505]=16'hc4ae;
aud[22506]=16'hc4a6;
aud[22507]=16'hc49e;
aud[22508]=16'hc496;
aud[22509]=16'hc48e;
aud[22510]=16'hc486;
aud[22511]=16'hc47f;
aud[22512]=16'hc477;
aud[22513]=16'hc46f;
aud[22514]=16'hc467;
aud[22515]=16'hc45f;
aud[22516]=16'hc457;
aud[22517]=16'hc450;
aud[22518]=16'hc448;
aud[22519]=16'hc440;
aud[22520]=16'hc439;
aud[22521]=16'hc431;
aud[22522]=16'hc429;
aud[22523]=16'hc422;
aud[22524]=16'hc41a;
aud[22525]=16'hc413;
aud[22526]=16'hc40b;
aud[22527]=16'hc404;
aud[22528]=16'hc3fc;
aud[22529]=16'hc3f5;
aud[22530]=16'hc3ed;
aud[22531]=16'hc3e6;
aud[22532]=16'hc3df;
aud[22533]=16'hc3d7;
aud[22534]=16'hc3d0;
aud[22535]=16'hc3c9;
aud[22536]=16'hc3c1;
aud[22537]=16'hc3ba;
aud[22538]=16'hc3b3;
aud[22539]=16'hc3ac;
aud[22540]=16'hc3a5;
aud[22541]=16'hc39d;
aud[22542]=16'hc396;
aud[22543]=16'hc38f;
aud[22544]=16'hc388;
aud[22545]=16'hc381;
aud[22546]=16'hc37a;
aud[22547]=16'hc373;
aud[22548]=16'hc36c;
aud[22549]=16'hc365;
aud[22550]=16'hc35f;
aud[22551]=16'hc358;
aud[22552]=16'hc351;
aud[22553]=16'hc34a;
aud[22554]=16'hc343;
aud[22555]=16'hc33d;
aud[22556]=16'hc336;
aud[22557]=16'hc32f;
aud[22558]=16'hc329;
aud[22559]=16'hc322;
aud[22560]=16'hc31b;
aud[22561]=16'hc315;
aud[22562]=16'hc30e;
aud[22563]=16'hc308;
aud[22564]=16'hc301;
aud[22565]=16'hc2fb;
aud[22566]=16'hc2f4;
aud[22567]=16'hc2ee;
aud[22568]=16'hc2e7;
aud[22569]=16'hc2e1;
aud[22570]=16'hc2db;
aud[22571]=16'hc2d4;
aud[22572]=16'hc2ce;
aud[22573]=16'hc2c8;
aud[22574]=16'hc2c1;
aud[22575]=16'hc2bb;
aud[22576]=16'hc2b5;
aud[22577]=16'hc2af;
aud[22578]=16'hc2a9;
aud[22579]=16'hc2a3;
aud[22580]=16'hc29d;
aud[22581]=16'hc297;
aud[22582]=16'hc291;
aud[22583]=16'hc28b;
aud[22584]=16'hc285;
aud[22585]=16'hc27f;
aud[22586]=16'hc279;
aud[22587]=16'hc273;
aud[22588]=16'hc26d;
aud[22589]=16'hc267;
aud[22590]=16'hc261;
aud[22591]=16'hc25c;
aud[22592]=16'hc256;
aud[22593]=16'hc250;
aud[22594]=16'hc24a;
aud[22595]=16'hc245;
aud[22596]=16'hc23f;
aud[22597]=16'hc239;
aud[22598]=16'hc234;
aud[22599]=16'hc22e;
aud[22600]=16'hc229;
aud[22601]=16'hc223;
aud[22602]=16'hc21e;
aud[22603]=16'hc218;
aud[22604]=16'hc213;
aud[22605]=16'hc20d;
aud[22606]=16'hc208;
aud[22607]=16'hc203;
aud[22608]=16'hc1fd;
aud[22609]=16'hc1f8;
aud[22610]=16'hc1f3;
aud[22611]=16'hc1ee;
aud[22612]=16'hc1e8;
aud[22613]=16'hc1e3;
aud[22614]=16'hc1de;
aud[22615]=16'hc1d9;
aud[22616]=16'hc1d4;
aud[22617]=16'hc1cf;
aud[22618]=16'hc1ca;
aud[22619]=16'hc1c5;
aud[22620]=16'hc1c0;
aud[22621]=16'hc1bb;
aud[22622]=16'hc1b6;
aud[22623]=16'hc1b1;
aud[22624]=16'hc1ac;
aud[22625]=16'hc1a7;
aud[22626]=16'hc1a2;
aud[22627]=16'hc19e;
aud[22628]=16'hc199;
aud[22629]=16'hc194;
aud[22630]=16'hc18f;
aud[22631]=16'hc18b;
aud[22632]=16'hc186;
aud[22633]=16'hc181;
aud[22634]=16'hc17d;
aud[22635]=16'hc178;
aud[22636]=16'hc174;
aud[22637]=16'hc16f;
aud[22638]=16'hc16b;
aud[22639]=16'hc166;
aud[22640]=16'hc162;
aud[22641]=16'hc15d;
aud[22642]=16'hc159;
aud[22643]=16'hc154;
aud[22644]=16'hc150;
aud[22645]=16'hc14c;
aud[22646]=16'hc147;
aud[22647]=16'hc143;
aud[22648]=16'hc13f;
aud[22649]=16'hc13b;
aud[22650]=16'hc137;
aud[22651]=16'hc133;
aud[22652]=16'hc12e;
aud[22653]=16'hc12a;
aud[22654]=16'hc126;
aud[22655]=16'hc122;
aud[22656]=16'hc11e;
aud[22657]=16'hc11a;
aud[22658]=16'hc116;
aud[22659]=16'hc112;
aud[22660]=16'hc10e;
aud[22661]=16'hc10b;
aud[22662]=16'hc107;
aud[22663]=16'hc103;
aud[22664]=16'hc0ff;
aud[22665]=16'hc0fb;
aud[22666]=16'hc0f8;
aud[22667]=16'hc0f4;
aud[22668]=16'hc0f0;
aud[22669]=16'hc0ed;
aud[22670]=16'hc0e9;
aud[22671]=16'hc0e5;
aud[22672]=16'hc0e2;
aud[22673]=16'hc0de;
aud[22674]=16'hc0db;
aud[22675]=16'hc0d7;
aud[22676]=16'hc0d4;
aud[22677]=16'hc0d0;
aud[22678]=16'hc0cd;
aud[22679]=16'hc0ca;
aud[22680]=16'hc0c6;
aud[22681]=16'hc0c3;
aud[22682]=16'hc0c0;
aud[22683]=16'hc0bd;
aud[22684]=16'hc0b9;
aud[22685]=16'hc0b6;
aud[22686]=16'hc0b3;
aud[22687]=16'hc0b0;
aud[22688]=16'hc0ad;
aud[22689]=16'hc0aa;
aud[22690]=16'hc0a6;
aud[22691]=16'hc0a3;
aud[22692]=16'hc0a0;
aud[22693]=16'hc09d;
aud[22694]=16'hc09b;
aud[22695]=16'hc098;
aud[22696]=16'hc095;
aud[22697]=16'hc092;
aud[22698]=16'hc08f;
aud[22699]=16'hc08c;
aud[22700]=16'hc089;
aud[22701]=16'hc087;
aud[22702]=16'hc084;
aud[22703]=16'hc081;
aud[22704]=16'hc07f;
aud[22705]=16'hc07c;
aud[22706]=16'hc079;
aud[22707]=16'hc077;
aud[22708]=16'hc074;
aud[22709]=16'hc072;
aud[22710]=16'hc06f;
aud[22711]=16'hc06d;
aud[22712]=16'hc06a;
aud[22713]=16'hc068;
aud[22714]=16'hc065;
aud[22715]=16'hc063;
aud[22716]=16'hc061;
aud[22717]=16'hc05e;
aud[22718]=16'hc05c;
aud[22719]=16'hc05a;
aud[22720]=16'hc058;
aud[22721]=16'hc055;
aud[22722]=16'hc053;
aud[22723]=16'hc051;
aud[22724]=16'hc04f;
aud[22725]=16'hc04d;
aud[22726]=16'hc04b;
aud[22727]=16'hc049;
aud[22728]=16'hc047;
aud[22729]=16'hc045;
aud[22730]=16'hc043;
aud[22731]=16'hc041;
aud[22732]=16'hc03f;
aud[22733]=16'hc03d;
aud[22734]=16'hc03b;
aud[22735]=16'hc039;
aud[22736]=16'hc038;
aud[22737]=16'hc036;
aud[22738]=16'hc034;
aud[22739]=16'hc033;
aud[22740]=16'hc031;
aud[22741]=16'hc02f;
aud[22742]=16'hc02e;
aud[22743]=16'hc02c;
aud[22744]=16'hc02a;
aud[22745]=16'hc029;
aud[22746]=16'hc027;
aud[22747]=16'hc026;
aud[22748]=16'hc024;
aud[22749]=16'hc023;
aud[22750]=16'hc022;
aud[22751]=16'hc020;
aud[22752]=16'hc01f;
aud[22753]=16'hc01e;
aud[22754]=16'hc01c;
aud[22755]=16'hc01b;
aud[22756]=16'hc01a;
aud[22757]=16'hc019;
aud[22758]=16'hc018;
aud[22759]=16'hc016;
aud[22760]=16'hc015;
aud[22761]=16'hc014;
aud[22762]=16'hc013;
aud[22763]=16'hc012;
aud[22764]=16'hc011;
aud[22765]=16'hc010;
aud[22766]=16'hc00f;
aud[22767]=16'hc00e;
aud[22768]=16'hc00d;
aud[22769]=16'hc00d;
aud[22770]=16'hc00c;
aud[22771]=16'hc00b;
aud[22772]=16'hc00a;
aud[22773]=16'hc009;
aud[22774]=16'hc009;
aud[22775]=16'hc008;
aud[22776]=16'hc007;
aud[22777]=16'hc007;
aud[22778]=16'hc006;
aud[22779]=16'hc006;
aud[22780]=16'hc005;
aud[22781]=16'hc005;
aud[22782]=16'hc004;
aud[22783]=16'hc004;
aud[22784]=16'hc003;
aud[22785]=16'hc003;
aud[22786]=16'hc002;
aud[22787]=16'hc002;
aud[22788]=16'hc002;
aud[22789]=16'hc001;
aud[22790]=16'hc001;
aud[22791]=16'hc001;
aud[22792]=16'hc001;
aud[22793]=16'hc001;
aud[22794]=16'hc000;
aud[22795]=16'hc000;
aud[22796]=16'hc000;
aud[22797]=16'hc000;
aud[22798]=16'hc000;
aud[22799]=16'hc000;
aud[22800]=16'hc000;
aud[22801]=16'hc000;
aud[22802]=16'hc000;
aud[22803]=16'hc000;
aud[22804]=16'hc000;
aud[22805]=16'hc001;
aud[22806]=16'hc001;
aud[22807]=16'hc001;
aud[22808]=16'hc001;
aud[22809]=16'hc001;
aud[22810]=16'hc002;
aud[22811]=16'hc002;
aud[22812]=16'hc002;
aud[22813]=16'hc003;
aud[22814]=16'hc003;
aud[22815]=16'hc004;
aud[22816]=16'hc004;
aud[22817]=16'hc005;
aud[22818]=16'hc005;
aud[22819]=16'hc006;
aud[22820]=16'hc006;
aud[22821]=16'hc007;
aud[22822]=16'hc007;
aud[22823]=16'hc008;
aud[22824]=16'hc009;
aud[22825]=16'hc009;
aud[22826]=16'hc00a;
aud[22827]=16'hc00b;
aud[22828]=16'hc00c;
aud[22829]=16'hc00d;
aud[22830]=16'hc00d;
aud[22831]=16'hc00e;
aud[22832]=16'hc00f;
aud[22833]=16'hc010;
aud[22834]=16'hc011;
aud[22835]=16'hc012;
aud[22836]=16'hc013;
aud[22837]=16'hc014;
aud[22838]=16'hc015;
aud[22839]=16'hc016;
aud[22840]=16'hc018;
aud[22841]=16'hc019;
aud[22842]=16'hc01a;
aud[22843]=16'hc01b;
aud[22844]=16'hc01c;
aud[22845]=16'hc01e;
aud[22846]=16'hc01f;
aud[22847]=16'hc020;
aud[22848]=16'hc022;
aud[22849]=16'hc023;
aud[22850]=16'hc024;
aud[22851]=16'hc026;
aud[22852]=16'hc027;
aud[22853]=16'hc029;
aud[22854]=16'hc02a;
aud[22855]=16'hc02c;
aud[22856]=16'hc02e;
aud[22857]=16'hc02f;
aud[22858]=16'hc031;
aud[22859]=16'hc033;
aud[22860]=16'hc034;
aud[22861]=16'hc036;
aud[22862]=16'hc038;
aud[22863]=16'hc039;
aud[22864]=16'hc03b;
aud[22865]=16'hc03d;
aud[22866]=16'hc03f;
aud[22867]=16'hc041;
aud[22868]=16'hc043;
aud[22869]=16'hc045;
aud[22870]=16'hc047;
aud[22871]=16'hc049;
aud[22872]=16'hc04b;
aud[22873]=16'hc04d;
aud[22874]=16'hc04f;
aud[22875]=16'hc051;
aud[22876]=16'hc053;
aud[22877]=16'hc055;
aud[22878]=16'hc058;
aud[22879]=16'hc05a;
aud[22880]=16'hc05c;
aud[22881]=16'hc05e;
aud[22882]=16'hc061;
aud[22883]=16'hc063;
aud[22884]=16'hc065;
aud[22885]=16'hc068;
aud[22886]=16'hc06a;
aud[22887]=16'hc06d;
aud[22888]=16'hc06f;
aud[22889]=16'hc072;
aud[22890]=16'hc074;
aud[22891]=16'hc077;
aud[22892]=16'hc079;
aud[22893]=16'hc07c;
aud[22894]=16'hc07f;
aud[22895]=16'hc081;
aud[22896]=16'hc084;
aud[22897]=16'hc087;
aud[22898]=16'hc089;
aud[22899]=16'hc08c;
aud[22900]=16'hc08f;
aud[22901]=16'hc092;
aud[22902]=16'hc095;
aud[22903]=16'hc098;
aud[22904]=16'hc09b;
aud[22905]=16'hc09d;
aud[22906]=16'hc0a0;
aud[22907]=16'hc0a3;
aud[22908]=16'hc0a6;
aud[22909]=16'hc0aa;
aud[22910]=16'hc0ad;
aud[22911]=16'hc0b0;
aud[22912]=16'hc0b3;
aud[22913]=16'hc0b6;
aud[22914]=16'hc0b9;
aud[22915]=16'hc0bd;
aud[22916]=16'hc0c0;
aud[22917]=16'hc0c3;
aud[22918]=16'hc0c6;
aud[22919]=16'hc0ca;
aud[22920]=16'hc0cd;
aud[22921]=16'hc0d0;
aud[22922]=16'hc0d4;
aud[22923]=16'hc0d7;
aud[22924]=16'hc0db;
aud[22925]=16'hc0de;
aud[22926]=16'hc0e2;
aud[22927]=16'hc0e5;
aud[22928]=16'hc0e9;
aud[22929]=16'hc0ed;
aud[22930]=16'hc0f0;
aud[22931]=16'hc0f4;
aud[22932]=16'hc0f8;
aud[22933]=16'hc0fb;
aud[22934]=16'hc0ff;
aud[22935]=16'hc103;
aud[22936]=16'hc107;
aud[22937]=16'hc10b;
aud[22938]=16'hc10e;
aud[22939]=16'hc112;
aud[22940]=16'hc116;
aud[22941]=16'hc11a;
aud[22942]=16'hc11e;
aud[22943]=16'hc122;
aud[22944]=16'hc126;
aud[22945]=16'hc12a;
aud[22946]=16'hc12e;
aud[22947]=16'hc133;
aud[22948]=16'hc137;
aud[22949]=16'hc13b;
aud[22950]=16'hc13f;
aud[22951]=16'hc143;
aud[22952]=16'hc147;
aud[22953]=16'hc14c;
aud[22954]=16'hc150;
aud[22955]=16'hc154;
aud[22956]=16'hc159;
aud[22957]=16'hc15d;
aud[22958]=16'hc162;
aud[22959]=16'hc166;
aud[22960]=16'hc16b;
aud[22961]=16'hc16f;
aud[22962]=16'hc174;
aud[22963]=16'hc178;
aud[22964]=16'hc17d;
aud[22965]=16'hc181;
aud[22966]=16'hc186;
aud[22967]=16'hc18b;
aud[22968]=16'hc18f;
aud[22969]=16'hc194;
aud[22970]=16'hc199;
aud[22971]=16'hc19e;
aud[22972]=16'hc1a2;
aud[22973]=16'hc1a7;
aud[22974]=16'hc1ac;
aud[22975]=16'hc1b1;
aud[22976]=16'hc1b6;
aud[22977]=16'hc1bb;
aud[22978]=16'hc1c0;
aud[22979]=16'hc1c5;
aud[22980]=16'hc1ca;
aud[22981]=16'hc1cf;
aud[22982]=16'hc1d4;
aud[22983]=16'hc1d9;
aud[22984]=16'hc1de;
aud[22985]=16'hc1e3;
aud[22986]=16'hc1e8;
aud[22987]=16'hc1ee;
aud[22988]=16'hc1f3;
aud[22989]=16'hc1f8;
aud[22990]=16'hc1fd;
aud[22991]=16'hc203;
aud[22992]=16'hc208;
aud[22993]=16'hc20d;
aud[22994]=16'hc213;
aud[22995]=16'hc218;
aud[22996]=16'hc21e;
aud[22997]=16'hc223;
aud[22998]=16'hc229;
aud[22999]=16'hc22e;
aud[23000]=16'hc234;
aud[23001]=16'hc239;
aud[23002]=16'hc23f;
aud[23003]=16'hc245;
aud[23004]=16'hc24a;
aud[23005]=16'hc250;
aud[23006]=16'hc256;
aud[23007]=16'hc25c;
aud[23008]=16'hc261;
aud[23009]=16'hc267;
aud[23010]=16'hc26d;
aud[23011]=16'hc273;
aud[23012]=16'hc279;
aud[23013]=16'hc27f;
aud[23014]=16'hc285;
aud[23015]=16'hc28b;
aud[23016]=16'hc291;
aud[23017]=16'hc297;
aud[23018]=16'hc29d;
aud[23019]=16'hc2a3;
aud[23020]=16'hc2a9;
aud[23021]=16'hc2af;
aud[23022]=16'hc2b5;
aud[23023]=16'hc2bb;
aud[23024]=16'hc2c1;
aud[23025]=16'hc2c8;
aud[23026]=16'hc2ce;
aud[23027]=16'hc2d4;
aud[23028]=16'hc2db;
aud[23029]=16'hc2e1;
aud[23030]=16'hc2e7;
aud[23031]=16'hc2ee;
aud[23032]=16'hc2f4;
aud[23033]=16'hc2fb;
aud[23034]=16'hc301;
aud[23035]=16'hc308;
aud[23036]=16'hc30e;
aud[23037]=16'hc315;
aud[23038]=16'hc31b;
aud[23039]=16'hc322;
aud[23040]=16'hc329;
aud[23041]=16'hc32f;
aud[23042]=16'hc336;
aud[23043]=16'hc33d;
aud[23044]=16'hc343;
aud[23045]=16'hc34a;
aud[23046]=16'hc351;
aud[23047]=16'hc358;
aud[23048]=16'hc35f;
aud[23049]=16'hc365;
aud[23050]=16'hc36c;
aud[23051]=16'hc373;
aud[23052]=16'hc37a;
aud[23053]=16'hc381;
aud[23054]=16'hc388;
aud[23055]=16'hc38f;
aud[23056]=16'hc396;
aud[23057]=16'hc39d;
aud[23058]=16'hc3a5;
aud[23059]=16'hc3ac;
aud[23060]=16'hc3b3;
aud[23061]=16'hc3ba;
aud[23062]=16'hc3c1;
aud[23063]=16'hc3c9;
aud[23064]=16'hc3d0;
aud[23065]=16'hc3d7;
aud[23066]=16'hc3df;
aud[23067]=16'hc3e6;
aud[23068]=16'hc3ed;
aud[23069]=16'hc3f5;
aud[23070]=16'hc3fc;
aud[23071]=16'hc404;
aud[23072]=16'hc40b;
aud[23073]=16'hc413;
aud[23074]=16'hc41a;
aud[23075]=16'hc422;
aud[23076]=16'hc429;
aud[23077]=16'hc431;
aud[23078]=16'hc439;
aud[23079]=16'hc440;
aud[23080]=16'hc448;
aud[23081]=16'hc450;
aud[23082]=16'hc457;
aud[23083]=16'hc45f;
aud[23084]=16'hc467;
aud[23085]=16'hc46f;
aud[23086]=16'hc477;
aud[23087]=16'hc47f;
aud[23088]=16'hc486;
aud[23089]=16'hc48e;
aud[23090]=16'hc496;
aud[23091]=16'hc49e;
aud[23092]=16'hc4a6;
aud[23093]=16'hc4ae;
aud[23094]=16'hc4b6;
aud[23095]=16'hc4bf;
aud[23096]=16'hc4c7;
aud[23097]=16'hc4cf;
aud[23098]=16'hc4d7;
aud[23099]=16'hc4df;
aud[23100]=16'hc4e7;
aud[23101]=16'hc4f0;
aud[23102]=16'hc4f8;
aud[23103]=16'hc500;
aud[23104]=16'hc509;
aud[23105]=16'hc511;
aud[23106]=16'hc519;
aud[23107]=16'hc522;
aud[23108]=16'hc52a;
aud[23109]=16'hc533;
aud[23110]=16'hc53b;
aud[23111]=16'hc544;
aud[23112]=16'hc54c;
aud[23113]=16'hc555;
aud[23114]=16'hc55d;
aud[23115]=16'hc566;
aud[23116]=16'hc56e;
aud[23117]=16'hc577;
aud[23118]=16'hc580;
aud[23119]=16'hc588;
aud[23120]=16'hc591;
aud[23121]=16'hc59a;
aud[23122]=16'hc5a3;
aud[23123]=16'hc5ac;
aud[23124]=16'hc5b4;
aud[23125]=16'hc5bd;
aud[23126]=16'hc5c6;
aud[23127]=16'hc5cf;
aud[23128]=16'hc5d8;
aud[23129]=16'hc5e1;
aud[23130]=16'hc5ea;
aud[23131]=16'hc5f3;
aud[23132]=16'hc5fc;
aud[23133]=16'hc605;
aud[23134]=16'hc60e;
aud[23135]=16'hc617;
aud[23136]=16'hc620;
aud[23137]=16'hc62a;
aud[23138]=16'hc633;
aud[23139]=16'hc63c;
aud[23140]=16'hc645;
aud[23141]=16'hc64f;
aud[23142]=16'hc658;
aud[23143]=16'hc661;
aud[23144]=16'hc66b;
aud[23145]=16'hc674;
aud[23146]=16'hc67d;
aud[23147]=16'hc687;
aud[23148]=16'hc690;
aud[23149]=16'hc69a;
aud[23150]=16'hc6a3;
aud[23151]=16'hc6ad;
aud[23152]=16'hc6b6;
aud[23153]=16'hc6c0;
aud[23154]=16'hc6c9;
aud[23155]=16'hc6d3;
aud[23156]=16'hc6dd;
aud[23157]=16'hc6e6;
aud[23158]=16'hc6f0;
aud[23159]=16'hc6fa;
aud[23160]=16'hc703;
aud[23161]=16'hc70d;
aud[23162]=16'hc717;
aud[23163]=16'hc721;
aud[23164]=16'hc72b;
aud[23165]=16'hc735;
aud[23166]=16'hc73f;
aud[23167]=16'hc748;
aud[23168]=16'hc752;
aud[23169]=16'hc75c;
aud[23170]=16'hc766;
aud[23171]=16'hc770;
aud[23172]=16'hc77a;
aud[23173]=16'hc785;
aud[23174]=16'hc78f;
aud[23175]=16'hc799;
aud[23176]=16'hc7a3;
aud[23177]=16'hc7ad;
aud[23178]=16'hc7b7;
aud[23179]=16'hc7c1;
aud[23180]=16'hc7cc;
aud[23181]=16'hc7d6;
aud[23182]=16'hc7e0;
aud[23183]=16'hc7eb;
aud[23184]=16'hc7f5;
aud[23185]=16'hc7ff;
aud[23186]=16'hc80a;
aud[23187]=16'hc814;
aud[23188]=16'hc81f;
aud[23189]=16'hc829;
aud[23190]=16'hc834;
aud[23191]=16'hc83e;
aud[23192]=16'hc849;
aud[23193]=16'hc853;
aud[23194]=16'hc85e;
aud[23195]=16'hc868;
aud[23196]=16'hc873;
aud[23197]=16'hc87e;
aud[23198]=16'hc888;
aud[23199]=16'hc893;
aud[23200]=16'hc89e;
aud[23201]=16'hc8a9;
aud[23202]=16'hc8b3;
aud[23203]=16'hc8be;
aud[23204]=16'hc8c9;
aud[23205]=16'hc8d4;
aud[23206]=16'hc8df;
aud[23207]=16'hc8ea;
aud[23208]=16'hc8f5;
aud[23209]=16'hc8ff;
aud[23210]=16'hc90a;
aud[23211]=16'hc915;
aud[23212]=16'hc920;
aud[23213]=16'hc92c;
aud[23214]=16'hc937;
aud[23215]=16'hc942;
aud[23216]=16'hc94d;
aud[23217]=16'hc958;
aud[23218]=16'hc963;
aud[23219]=16'hc96e;
aud[23220]=16'hc97a;
aud[23221]=16'hc985;
aud[23222]=16'hc990;
aud[23223]=16'hc99b;
aud[23224]=16'hc9a7;
aud[23225]=16'hc9b2;
aud[23226]=16'hc9bd;
aud[23227]=16'hc9c9;
aud[23228]=16'hc9d4;
aud[23229]=16'hc9e0;
aud[23230]=16'hc9eb;
aud[23231]=16'hc9f7;
aud[23232]=16'hca02;
aud[23233]=16'hca0e;
aud[23234]=16'hca19;
aud[23235]=16'hca25;
aud[23236]=16'hca30;
aud[23237]=16'hca3c;
aud[23238]=16'hca48;
aud[23239]=16'hca53;
aud[23240]=16'hca5f;
aud[23241]=16'hca6b;
aud[23242]=16'hca76;
aud[23243]=16'hca82;
aud[23244]=16'hca8e;
aud[23245]=16'hca9a;
aud[23246]=16'hcaa6;
aud[23247]=16'hcab1;
aud[23248]=16'hcabd;
aud[23249]=16'hcac9;
aud[23250]=16'hcad5;
aud[23251]=16'hcae1;
aud[23252]=16'hcaed;
aud[23253]=16'hcaf9;
aud[23254]=16'hcb05;
aud[23255]=16'hcb11;
aud[23256]=16'hcb1d;
aud[23257]=16'hcb29;
aud[23258]=16'hcb35;
aud[23259]=16'hcb42;
aud[23260]=16'hcb4e;
aud[23261]=16'hcb5a;
aud[23262]=16'hcb66;
aud[23263]=16'hcb72;
aud[23264]=16'hcb7f;
aud[23265]=16'hcb8b;
aud[23266]=16'hcb97;
aud[23267]=16'hcba3;
aud[23268]=16'hcbb0;
aud[23269]=16'hcbbc;
aud[23270]=16'hcbc9;
aud[23271]=16'hcbd5;
aud[23272]=16'hcbe1;
aud[23273]=16'hcbee;
aud[23274]=16'hcbfa;
aud[23275]=16'hcc07;
aud[23276]=16'hcc13;
aud[23277]=16'hcc20;
aud[23278]=16'hcc2c;
aud[23279]=16'hcc39;
aud[23280]=16'hcc46;
aud[23281]=16'hcc52;
aud[23282]=16'hcc5f;
aud[23283]=16'hcc6c;
aud[23284]=16'hcc78;
aud[23285]=16'hcc85;
aud[23286]=16'hcc92;
aud[23287]=16'hcc9f;
aud[23288]=16'hccab;
aud[23289]=16'hccb8;
aud[23290]=16'hccc5;
aud[23291]=16'hccd2;
aud[23292]=16'hccdf;
aud[23293]=16'hccec;
aud[23294]=16'hccf9;
aud[23295]=16'hcd06;
aud[23296]=16'hcd13;
aud[23297]=16'hcd20;
aud[23298]=16'hcd2d;
aud[23299]=16'hcd3a;
aud[23300]=16'hcd47;
aud[23301]=16'hcd54;
aud[23302]=16'hcd61;
aud[23303]=16'hcd6e;
aud[23304]=16'hcd7b;
aud[23305]=16'hcd88;
aud[23306]=16'hcd96;
aud[23307]=16'hcda3;
aud[23308]=16'hcdb0;
aud[23309]=16'hcdbd;
aud[23310]=16'hcdcb;
aud[23311]=16'hcdd8;
aud[23312]=16'hcde5;
aud[23313]=16'hcdf3;
aud[23314]=16'hce00;
aud[23315]=16'hce0d;
aud[23316]=16'hce1b;
aud[23317]=16'hce28;
aud[23318]=16'hce36;
aud[23319]=16'hce43;
aud[23320]=16'hce51;
aud[23321]=16'hce5e;
aud[23322]=16'hce6c;
aud[23323]=16'hce79;
aud[23324]=16'hce87;
aud[23325]=16'hce95;
aud[23326]=16'hcea2;
aud[23327]=16'hceb0;
aud[23328]=16'hcebe;
aud[23329]=16'hcecb;
aud[23330]=16'hced9;
aud[23331]=16'hcee7;
aud[23332]=16'hcef5;
aud[23333]=16'hcf02;
aud[23334]=16'hcf10;
aud[23335]=16'hcf1e;
aud[23336]=16'hcf2c;
aud[23337]=16'hcf3a;
aud[23338]=16'hcf48;
aud[23339]=16'hcf56;
aud[23340]=16'hcf63;
aud[23341]=16'hcf71;
aud[23342]=16'hcf7f;
aud[23343]=16'hcf8d;
aud[23344]=16'hcf9b;
aud[23345]=16'hcfa9;
aud[23346]=16'hcfb8;
aud[23347]=16'hcfc6;
aud[23348]=16'hcfd4;
aud[23349]=16'hcfe2;
aud[23350]=16'hcff0;
aud[23351]=16'hcffe;
aud[23352]=16'hd00c;
aud[23353]=16'hd01b;
aud[23354]=16'hd029;
aud[23355]=16'hd037;
aud[23356]=16'hd045;
aud[23357]=16'hd054;
aud[23358]=16'hd062;
aud[23359]=16'hd070;
aud[23360]=16'hd07f;
aud[23361]=16'hd08d;
aud[23362]=16'hd09b;
aud[23363]=16'hd0aa;
aud[23364]=16'hd0b8;
aud[23365]=16'hd0c7;
aud[23366]=16'hd0d5;
aud[23367]=16'hd0e4;
aud[23368]=16'hd0f2;
aud[23369]=16'hd101;
aud[23370]=16'hd10f;
aud[23371]=16'hd11e;
aud[23372]=16'hd12d;
aud[23373]=16'hd13b;
aud[23374]=16'hd14a;
aud[23375]=16'hd159;
aud[23376]=16'hd167;
aud[23377]=16'hd176;
aud[23378]=16'hd185;
aud[23379]=16'hd193;
aud[23380]=16'hd1a2;
aud[23381]=16'hd1b1;
aud[23382]=16'hd1c0;
aud[23383]=16'hd1cf;
aud[23384]=16'hd1de;
aud[23385]=16'hd1ec;
aud[23386]=16'hd1fb;
aud[23387]=16'hd20a;
aud[23388]=16'hd219;
aud[23389]=16'hd228;
aud[23390]=16'hd237;
aud[23391]=16'hd246;
aud[23392]=16'hd255;
aud[23393]=16'hd264;
aud[23394]=16'hd273;
aud[23395]=16'hd282;
aud[23396]=16'hd291;
aud[23397]=16'hd2a0;
aud[23398]=16'hd2b0;
aud[23399]=16'hd2bf;
aud[23400]=16'hd2ce;
aud[23401]=16'hd2dd;
aud[23402]=16'hd2ec;
aud[23403]=16'hd2fc;
aud[23404]=16'hd30b;
aud[23405]=16'hd31a;
aud[23406]=16'hd329;
aud[23407]=16'hd339;
aud[23408]=16'hd348;
aud[23409]=16'hd357;
aud[23410]=16'hd367;
aud[23411]=16'hd376;
aud[23412]=16'hd386;
aud[23413]=16'hd395;
aud[23414]=16'hd3a4;
aud[23415]=16'hd3b4;
aud[23416]=16'hd3c3;
aud[23417]=16'hd3d3;
aud[23418]=16'hd3e2;
aud[23419]=16'hd3f2;
aud[23420]=16'hd402;
aud[23421]=16'hd411;
aud[23422]=16'hd421;
aud[23423]=16'hd430;
aud[23424]=16'hd440;
aud[23425]=16'hd450;
aud[23426]=16'hd45f;
aud[23427]=16'hd46f;
aud[23428]=16'hd47f;
aud[23429]=16'hd48f;
aud[23430]=16'hd49e;
aud[23431]=16'hd4ae;
aud[23432]=16'hd4be;
aud[23433]=16'hd4ce;
aud[23434]=16'hd4de;
aud[23435]=16'hd4ed;
aud[23436]=16'hd4fd;
aud[23437]=16'hd50d;
aud[23438]=16'hd51d;
aud[23439]=16'hd52d;
aud[23440]=16'hd53d;
aud[23441]=16'hd54d;
aud[23442]=16'hd55d;
aud[23443]=16'hd56d;
aud[23444]=16'hd57d;
aud[23445]=16'hd58d;
aud[23446]=16'hd59d;
aud[23447]=16'hd5ad;
aud[23448]=16'hd5bd;
aud[23449]=16'hd5cd;
aud[23450]=16'hd5dd;
aud[23451]=16'hd5ee;
aud[23452]=16'hd5fe;
aud[23453]=16'hd60e;
aud[23454]=16'hd61e;
aud[23455]=16'hd62e;
aud[23456]=16'hd63f;
aud[23457]=16'hd64f;
aud[23458]=16'hd65f;
aud[23459]=16'hd66f;
aud[23460]=16'hd680;
aud[23461]=16'hd690;
aud[23462]=16'hd6a0;
aud[23463]=16'hd6b1;
aud[23464]=16'hd6c1;
aud[23465]=16'hd6d2;
aud[23466]=16'hd6e2;
aud[23467]=16'hd6f2;
aud[23468]=16'hd703;
aud[23469]=16'hd713;
aud[23470]=16'hd724;
aud[23471]=16'hd734;
aud[23472]=16'hd745;
aud[23473]=16'hd756;
aud[23474]=16'hd766;
aud[23475]=16'hd777;
aud[23476]=16'hd787;
aud[23477]=16'hd798;
aud[23478]=16'hd7a9;
aud[23479]=16'hd7b9;
aud[23480]=16'hd7ca;
aud[23481]=16'hd7db;
aud[23482]=16'hd7eb;
aud[23483]=16'hd7fc;
aud[23484]=16'hd80d;
aud[23485]=16'hd81e;
aud[23486]=16'hd82e;
aud[23487]=16'hd83f;
aud[23488]=16'hd850;
aud[23489]=16'hd861;
aud[23490]=16'hd872;
aud[23491]=16'hd882;
aud[23492]=16'hd893;
aud[23493]=16'hd8a4;
aud[23494]=16'hd8b5;
aud[23495]=16'hd8c6;
aud[23496]=16'hd8d7;
aud[23497]=16'hd8e8;
aud[23498]=16'hd8f9;
aud[23499]=16'hd90a;
aud[23500]=16'hd91b;
aud[23501]=16'hd92c;
aud[23502]=16'hd93d;
aud[23503]=16'hd94e;
aud[23504]=16'hd95f;
aud[23505]=16'hd970;
aud[23506]=16'hd982;
aud[23507]=16'hd993;
aud[23508]=16'hd9a4;
aud[23509]=16'hd9b5;
aud[23510]=16'hd9c6;
aud[23511]=16'hd9d7;
aud[23512]=16'hd9e9;
aud[23513]=16'hd9fa;
aud[23514]=16'hda0b;
aud[23515]=16'hda1c;
aud[23516]=16'hda2e;
aud[23517]=16'hda3f;
aud[23518]=16'hda50;
aud[23519]=16'hda62;
aud[23520]=16'hda73;
aud[23521]=16'hda84;
aud[23522]=16'hda96;
aud[23523]=16'hdaa7;
aud[23524]=16'hdab9;
aud[23525]=16'hdaca;
aud[23526]=16'hdadc;
aud[23527]=16'hdaed;
aud[23528]=16'hdaff;
aud[23529]=16'hdb10;
aud[23530]=16'hdb22;
aud[23531]=16'hdb33;
aud[23532]=16'hdb45;
aud[23533]=16'hdb56;
aud[23534]=16'hdb68;
aud[23535]=16'hdb79;
aud[23536]=16'hdb8b;
aud[23537]=16'hdb9d;
aud[23538]=16'hdbae;
aud[23539]=16'hdbc0;
aud[23540]=16'hdbd2;
aud[23541]=16'hdbe3;
aud[23542]=16'hdbf5;
aud[23543]=16'hdc07;
aud[23544]=16'hdc19;
aud[23545]=16'hdc2a;
aud[23546]=16'hdc3c;
aud[23547]=16'hdc4e;
aud[23548]=16'hdc60;
aud[23549]=16'hdc72;
aud[23550]=16'hdc83;
aud[23551]=16'hdc95;
aud[23552]=16'hdca7;
aud[23553]=16'hdcb9;
aud[23554]=16'hdccb;
aud[23555]=16'hdcdd;
aud[23556]=16'hdcef;
aud[23557]=16'hdd01;
aud[23558]=16'hdd13;
aud[23559]=16'hdd25;
aud[23560]=16'hdd37;
aud[23561]=16'hdd49;
aud[23562]=16'hdd5b;
aud[23563]=16'hdd6d;
aud[23564]=16'hdd7f;
aud[23565]=16'hdd91;
aud[23566]=16'hdda3;
aud[23567]=16'hddb5;
aud[23568]=16'hddc7;
aud[23569]=16'hddd9;
aud[23570]=16'hddeb;
aud[23571]=16'hddfe;
aud[23572]=16'hde10;
aud[23573]=16'hde22;
aud[23574]=16'hde34;
aud[23575]=16'hde46;
aud[23576]=16'hde59;
aud[23577]=16'hde6b;
aud[23578]=16'hde7d;
aud[23579]=16'hde8f;
aud[23580]=16'hdea2;
aud[23581]=16'hdeb4;
aud[23582]=16'hdec6;
aud[23583]=16'hded9;
aud[23584]=16'hdeeb;
aud[23585]=16'hdefd;
aud[23586]=16'hdf10;
aud[23587]=16'hdf22;
aud[23588]=16'hdf35;
aud[23589]=16'hdf47;
aud[23590]=16'hdf59;
aud[23591]=16'hdf6c;
aud[23592]=16'hdf7e;
aud[23593]=16'hdf91;
aud[23594]=16'hdfa3;
aud[23595]=16'hdfb6;
aud[23596]=16'hdfc8;
aud[23597]=16'hdfdb;
aud[23598]=16'hdfed;
aud[23599]=16'he000;
aud[23600]=16'he013;
aud[23601]=16'he025;
aud[23602]=16'he038;
aud[23603]=16'he04a;
aud[23604]=16'he05d;
aud[23605]=16'he070;
aud[23606]=16'he082;
aud[23607]=16'he095;
aud[23608]=16'he0a8;
aud[23609]=16'he0ba;
aud[23610]=16'he0cd;
aud[23611]=16'he0e0;
aud[23612]=16'he0f3;
aud[23613]=16'he105;
aud[23614]=16'he118;
aud[23615]=16'he12b;
aud[23616]=16'he13e;
aud[23617]=16'he151;
aud[23618]=16'he163;
aud[23619]=16'he176;
aud[23620]=16'he189;
aud[23621]=16'he19c;
aud[23622]=16'he1af;
aud[23623]=16'he1c2;
aud[23624]=16'he1d5;
aud[23625]=16'he1e8;
aud[23626]=16'he1fa;
aud[23627]=16'he20d;
aud[23628]=16'he220;
aud[23629]=16'he233;
aud[23630]=16'he246;
aud[23631]=16'he259;
aud[23632]=16'he26c;
aud[23633]=16'he27f;
aud[23634]=16'he292;
aud[23635]=16'he2a5;
aud[23636]=16'he2b9;
aud[23637]=16'he2cc;
aud[23638]=16'he2df;
aud[23639]=16'he2f2;
aud[23640]=16'he305;
aud[23641]=16'he318;
aud[23642]=16'he32b;
aud[23643]=16'he33e;
aud[23644]=16'he352;
aud[23645]=16'he365;
aud[23646]=16'he378;
aud[23647]=16'he38b;
aud[23648]=16'he39e;
aud[23649]=16'he3b2;
aud[23650]=16'he3c5;
aud[23651]=16'he3d8;
aud[23652]=16'he3eb;
aud[23653]=16'he3ff;
aud[23654]=16'he412;
aud[23655]=16'he425;
aud[23656]=16'he438;
aud[23657]=16'he44c;
aud[23658]=16'he45f;
aud[23659]=16'he473;
aud[23660]=16'he486;
aud[23661]=16'he499;
aud[23662]=16'he4ad;
aud[23663]=16'he4c0;
aud[23664]=16'he4d3;
aud[23665]=16'he4e7;
aud[23666]=16'he4fa;
aud[23667]=16'he50e;
aud[23668]=16'he521;
aud[23669]=16'he535;
aud[23670]=16'he548;
aud[23671]=16'he55c;
aud[23672]=16'he56f;
aud[23673]=16'he583;
aud[23674]=16'he596;
aud[23675]=16'he5aa;
aud[23676]=16'he5bd;
aud[23677]=16'he5d1;
aud[23678]=16'he5e4;
aud[23679]=16'he5f8;
aud[23680]=16'he60c;
aud[23681]=16'he61f;
aud[23682]=16'he633;
aud[23683]=16'he646;
aud[23684]=16'he65a;
aud[23685]=16'he66e;
aud[23686]=16'he681;
aud[23687]=16'he695;
aud[23688]=16'he6a9;
aud[23689]=16'he6bd;
aud[23690]=16'he6d0;
aud[23691]=16'he6e4;
aud[23692]=16'he6f8;
aud[23693]=16'he70b;
aud[23694]=16'he71f;
aud[23695]=16'he733;
aud[23696]=16'he747;
aud[23697]=16'he75b;
aud[23698]=16'he76e;
aud[23699]=16'he782;
aud[23700]=16'he796;
aud[23701]=16'he7aa;
aud[23702]=16'he7be;
aud[23703]=16'he7d1;
aud[23704]=16'he7e5;
aud[23705]=16'he7f9;
aud[23706]=16'he80d;
aud[23707]=16'he821;
aud[23708]=16'he835;
aud[23709]=16'he849;
aud[23710]=16'he85d;
aud[23711]=16'he871;
aud[23712]=16'he885;
aud[23713]=16'he899;
aud[23714]=16'he8ad;
aud[23715]=16'he8c0;
aud[23716]=16'he8d4;
aud[23717]=16'he8e8;
aud[23718]=16'he8fc;
aud[23719]=16'he910;
aud[23720]=16'he925;
aud[23721]=16'he939;
aud[23722]=16'he94d;
aud[23723]=16'he961;
aud[23724]=16'he975;
aud[23725]=16'he989;
aud[23726]=16'he99d;
aud[23727]=16'he9b1;
aud[23728]=16'he9c5;
aud[23729]=16'he9d9;
aud[23730]=16'he9ed;
aud[23731]=16'hea01;
aud[23732]=16'hea16;
aud[23733]=16'hea2a;
aud[23734]=16'hea3e;
aud[23735]=16'hea52;
aud[23736]=16'hea66;
aud[23737]=16'hea7a;
aud[23738]=16'hea8f;
aud[23739]=16'heaa3;
aud[23740]=16'heab7;
aud[23741]=16'heacb;
aud[23742]=16'heae0;
aud[23743]=16'heaf4;
aud[23744]=16'heb08;
aud[23745]=16'heb1c;
aud[23746]=16'heb31;
aud[23747]=16'heb45;
aud[23748]=16'heb59;
aud[23749]=16'heb6e;
aud[23750]=16'heb82;
aud[23751]=16'heb96;
aud[23752]=16'hebab;
aud[23753]=16'hebbf;
aud[23754]=16'hebd3;
aud[23755]=16'hebe8;
aud[23756]=16'hebfc;
aud[23757]=16'hec10;
aud[23758]=16'hec25;
aud[23759]=16'hec39;
aud[23760]=16'hec4d;
aud[23761]=16'hec62;
aud[23762]=16'hec76;
aud[23763]=16'hec8b;
aud[23764]=16'hec9f;
aud[23765]=16'hecb4;
aud[23766]=16'hecc8;
aud[23767]=16'hecdd;
aud[23768]=16'hecf1;
aud[23769]=16'hed05;
aud[23770]=16'hed1a;
aud[23771]=16'hed2e;
aud[23772]=16'hed43;
aud[23773]=16'hed57;
aud[23774]=16'hed6c;
aud[23775]=16'hed81;
aud[23776]=16'hed95;
aud[23777]=16'hedaa;
aud[23778]=16'hedbe;
aud[23779]=16'hedd3;
aud[23780]=16'hede7;
aud[23781]=16'hedfc;
aud[23782]=16'hee10;
aud[23783]=16'hee25;
aud[23784]=16'hee3a;
aud[23785]=16'hee4e;
aud[23786]=16'hee63;
aud[23787]=16'hee77;
aud[23788]=16'hee8c;
aud[23789]=16'heea1;
aud[23790]=16'heeb5;
aud[23791]=16'heeca;
aud[23792]=16'heedf;
aud[23793]=16'heef3;
aud[23794]=16'hef08;
aud[23795]=16'hef1d;
aud[23796]=16'hef31;
aud[23797]=16'hef46;
aud[23798]=16'hef5b;
aud[23799]=16'hef70;
aud[23800]=16'hef84;
aud[23801]=16'hef99;
aud[23802]=16'hefae;
aud[23803]=16'hefc2;
aud[23804]=16'hefd7;
aud[23805]=16'hefec;
aud[23806]=16'hf001;
aud[23807]=16'hf015;
aud[23808]=16'hf02a;
aud[23809]=16'hf03f;
aud[23810]=16'hf054;
aud[23811]=16'hf069;
aud[23812]=16'hf07d;
aud[23813]=16'hf092;
aud[23814]=16'hf0a7;
aud[23815]=16'hf0bc;
aud[23816]=16'hf0d1;
aud[23817]=16'hf0e6;
aud[23818]=16'hf0fa;
aud[23819]=16'hf10f;
aud[23820]=16'hf124;
aud[23821]=16'hf139;
aud[23822]=16'hf14e;
aud[23823]=16'hf163;
aud[23824]=16'hf178;
aud[23825]=16'hf18c;
aud[23826]=16'hf1a1;
aud[23827]=16'hf1b6;
aud[23828]=16'hf1cb;
aud[23829]=16'hf1e0;
aud[23830]=16'hf1f5;
aud[23831]=16'hf20a;
aud[23832]=16'hf21f;
aud[23833]=16'hf234;
aud[23834]=16'hf249;
aud[23835]=16'hf25e;
aud[23836]=16'hf273;
aud[23837]=16'hf288;
aud[23838]=16'hf29d;
aud[23839]=16'hf2b2;
aud[23840]=16'hf2c7;
aud[23841]=16'hf2dc;
aud[23842]=16'hf2f1;
aud[23843]=16'hf306;
aud[23844]=16'hf31b;
aud[23845]=16'hf330;
aud[23846]=16'hf345;
aud[23847]=16'hf35a;
aud[23848]=16'hf36f;
aud[23849]=16'hf384;
aud[23850]=16'hf399;
aud[23851]=16'hf3ae;
aud[23852]=16'hf3c3;
aud[23853]=16'hf3d8;
aud[23854]=16'hf3ed;
aud[23855]=16'hf402;
aud[23856]=16'hf417;
aud[23857]=16'hf42c;
aud[23858]=16'hf441;
aud[23859]=16'hf456;
aud[23860]=16'hf46b;
aud[23861]=16'hf480;
aud[23862]=16'hf496;
aud[23863]=16'hf4ab;
aud[23864]=16'hf4c0;
aud[23865]=16'hf4d5;
aud[23866]=16'hf4ea;
aud[23867]=16'hf4ff;
aud[23868]=16'hf514;
aud[23869]=16'hf529;
aud[23870]=16'hf53f;
aud[23871]=16'hf554;
aud[23872]=16'hf569;
aud[23873]=16'hf57e;
aud[23874]=16'hf593;
aud[23875]=16'hf5a8;
aud[23876]=16'hf5bd;
aud[23877]=16'hf5d3;
aud[23878]=16'hf5e8;
aud[23879]=16'hf5fd;
aud[23880]=16'hf612;
aud[23881]=16'hf627;
aud[23882]=16'hf63d;
aud[23883]=16'hf652;
aud[23884]=16'hf667;
aud[23885]=16'hf67c;
aud[23886]=16'hf691;
aud[23887]=16'hf6a7;
aud[23888]=16'hf6bc;
aud[23889]=16'hf6d1;
aud[23890]=16'hf6e6;
aud[23891]=16'hf6fb;
aud[23892]=16'hf711;
aud[23893]=16'hf726;
aud[23894]=16'hf73b;
aud[23895]=16'hf750;
aud[23896]=16'hf766;
aud[23897]=16'hf77b;
aud[23898]=16'hf790;
aud[23899]=16'hf7a5;
aud[23900]=16'hf7bb;
aud[23901]=16'hf7d0;
aud[23902]=16'hf7e5;
aud[23903]=16'hf7fb;
aud[23904]=16'hf810;
aud[23905]=16'hf825;
aud[23906]=16'hf83a;
aud[23907]=16'hf850;
aud[23908]=16'hf865;
aud[23909]=16'hf87a;
aud[23910]=16'hf890;
aud[23911]=16'hf8a5;
aud[23912]=16'hf8ba;
aud[23913]=16'hf8cf;
aud[23914]=16'hf8e5;
aud[23915]=16'hf8fa;
aud[23916]=16'hf90f;
aud[23917]=16'hf925;
aud[23918]=16'hf93a;
aud[23919]=16'hf94f;
aud[23920]=16'hf965;
aud[23921]=16'hf97a;
aud[23922]=16'hf98f;
aud[23923]=16'hf9a5;
aud[23924]=16'hf9ba;
aud[23925]=16'hf9cf;
aud[23926]=16'hf9e5;
aud[23927]=16'hf9fa;
aud[23928]=16'hfa0f;
aud[23929]=16'hfa25;
aud[23930]=16'hfa3a;
aud[23931]=16'hfa50;
aud[23932]=16'hfa65;
aud[23933]=16'hfa7a;
aud[23934]=16'hfa90;
aud[23935]=16'hfaa5;
aud[23936]=16'hfaba;
aud[23937]=16'hfad0;
aud[23938]=16'hfae5;
aud[23939]=16'hfafb;
aud[23940]=16'hfb10;
aud[23941]=16'hfb25;
aud[23942]=16'hfb3b;
aud[23943]=16'hfb50;
aud[23944]=16'hfb65;
aud[23945]=16'hfb7b;
aud[23946]=16'hfb90;
aud[23947]=16'hfba6;
aud[23948]=16'hfbbb;
aud[23949]=16'hfbd0;
aud[23950]=16'hfbe6;
aud[23951]=16'hfbfb;
aud[23952]=16'hfc11;
aud[23953]=16'hfc26;
aud[23954]=16'hfc3b;
aud[23955]=16'hfc51;
aud[23956]=16'hfc66;
aud[23957]=16'hfc7c;
aud[23958]=16'hfc91;
aud[23959]=16'hfca7;
aud[23960]=16'hfcbc;
aud[23961]=16'hfcd1;
aud[23962]=16'hfce7;
aud[23963]=16'hfcfc;
aud[23964]=16'hfd12;
aud[23965]=16'hfd27;
aud[23966]=16'hfd3c;
aud[23967]=16'hfd52;
aud[23968]=16'hfd67;
aud[23969]=16'hfd7d;
aud[23970]=16'hfd92;
aud[23971]=16'hfda8;
aud[23972]=16'hfdbd;
aud[23973]=16'hfdd2;
aud[23974]=16'hfde8;
aud[23975]=16'hfdfd;
aud[23976]=16'hfe13;
aud[23977]=16'hfe28;
aud[23978]=16'hfe3e;
aud[23979]=16'hfe53;
aud[23980]=16'hfe69;
aud[23981]=16'hfe7e;
aud[23982]=16'hfe93;
aud[23983]=16'hfea9;
aud[23984]=16'hfebe;
aud[23985]=16'hfed4;
aud[23986]=16'hfee9;
aud[23987]=16'hfeff;
aud[23988]=16'hff14;
aud[23989]=16'hff2a;
aud[23990]=16'hff3f;
aud[23991]=16'hff54;
aud[23992]=16'hff6a;
aud[23993]=16'hff7f;
aud[23994]=16'hff95;
aud[23995]=16'hffaa;
aud[23996]=16'hffc0;
aud[23997]=16'hffd5;
aud[23998]=16'hffeb;
aud[23999]=16'h0;
aud[24000]=16'h15;
aud[24001]=16'h2b;
aud[24002]=16'h40;
aud[24003]=16'h56;
aud[24004]=16'h6b;
aud[24005]=16'h81;
aud[24006]=16'h96;
aud[24007]=16'hac;
aud[24008]=16'hc1;
aud[24009]=16'hd6;
aud[24010]=16'hec;
aud[24011]=16'h101;
aud[24012]=16'h117;
aud[24013]=16'h12c;
aud[24014]=16'h142;
aud[24015]=16'h157;
aud[24016]=16'h16d;
aud[24017]=16'h182;
aud[24018]=16'h197;
aud[24019]=16'h1ad;
aud[24020]=16'h1c2;
aud[24021]=16'h1d8;
aud[24022]=16'h1ed;
aud[24023]=16'h203;
aud[24024]=16'h218;
aud[24025]=16'h22e;
aud[24026]=16'h243;
aud[24027]=16'h258;
aud[24028]=16'h26e;
aud[24029]=16'h283;
aud[24030]=16'h299;
aud[24031]=16'h2ae;
aud[24032]=16'h2c4;
aud[24033]=16'h2d9;
aud[24034]=16'h2ee;
aud[24035]=16'h304;
aud[24036]=16'h319;
aud[24037]=16'h32f;
aud[24038]=16'h344;
aud[24039]=16'h359;
aud[24040]=16'h36f;
aud[24041]=16'h384;
aud[24042]=16'h39a;
aud[24043]=16'h3af;
aud[24044]=16'h3c5;
aud[24045]=16'h3da;
aud[24046]=16'h3ef;
aud[24047]=16'h405;
aud[24048]=16'h41a;
aud[24049]=16'h430;
aud[24050]=16'h445;
aud[24051]=16'h45a;
aud[24052]=16'h470;
aud[24053]=16'h485;
aud[24054]=16'h49b;
aud[24055]=16'h4b0;
aud[24056]=16'h4c5;
aud[24057]=16'h4db;
aud[24058]=16'h4f0;
aud[24059]=16'h505;
aud[24060]=16'h51b;
aud[24061]=16'h530;
aud[24062]=16'h546;
aud[24063]=16'h55b;
aud[24064]=16'h570;
aud[24065]=16'h586;
aud[24066]=16'h59b;
aud[24067]=16'h5b0;
aud[24068]=16'h5c6;
aud[24069]=16'h5db;
aud[24070]=16'h5f1;
aud[24071]=16'h606;
aud[24072]=16'h61b;
aud[24073]=16'h631;
aud[24074]=16'h646;
aud[24075]=16'h65b;
aud[24076]=16'h671;
aud[24077]=16'h686;
aud[24078]=16'h69b;
aud[24079]=16'h6b1;
aud[24080]=16'h6c6;
aud[24081]=16'h6db;
aud[24082]=16'h6f1;
aud[24083]=16'h706;
aud[24084]=16'h71b;
aud[24085]=16'h731;
aud[24086]=16'h746;
aud[24087]=16'h75b;
aud[24088]=16'h770;
aud[24089]=16'h786;
aud[24090]=16'h79b;
aud[24091]=16'h7b0;
aud[24092]=16'h7c6;
aud[24093]=16'h7db;
aud[24094]=16'h7f0;
aud[24095]=16'h805;
aud[24096]=16'h81b;
aud[24097]=16'h830;
aud[24098]=16'h845;
aud[24099]=16'h85b;
aud[24100]=16'h870;
aud[24101]=16'h885;
aud[24102]=16'h89a;
aud[24103]=16'h8b0;
aud[24104]=16'h8c5;
aud[24105]=16'h8da;
aud[24106]=16'h8ef;
aud[24107]=16'h905;
aud[24108]=16'h91a;
aud[24109]=16'h92f;
aud[24110]=16'h944;
aud[24111]=16'h959;
aud[24112]=16'h96f;
aud[24113]=16'h984;
aud[24114]=16'h999;
aud[24115]=16'h9ae;
aud[24116]=16'h9c3;
aud[24117]=16'h9d9;
aud[24118]=16'h9ee;
aud[24119]=16'ha03;
aud[24120]=16'ha18;
aud[24121]=16'ha2d;
aud[24122]=16'ha43;
aud[24123]=16'ha58;
aud[24124]=16'ha6d;
aud[24125]=16'ha82;
aud[24126]=16'ha97;
aud[24127]=16'haac;
aud[24128]=16'hac1;
aud[24129]=16'had7;
aud[24130]=16'haec;
aud[24131]=16'hb01;
aud[24132]=16'hb16;
aud[24133]=16'hb2b;
aud[24134]=16'hb40;
aud[24135]=16'hb55;
aud[24136]=16'hb6a;
aud[24137]=16'hb80;
aud[24138]=16'hb95;
aud[24139]=16'hbaa;
aud[24140]=16'hbbf;
aud[24141]=16'hbd4;
aud[24142]=16'hbe9;
aud[24143]=16'hbfe;
aud[24144]=16'hc13;
aud[24145]=16'hc28;
aud[24146]=16'hc3d;
aud[24147]=16'hc52;
aud[24148]=16'hc67;
aud[24149]=16'hc7c;
aud[24150]=16'hc91;
aud[24151]=16'hca6;
aud[24152]=16'hcbb;
aud[24153]=16'hcd0;
aud[24154]=16'hce5;
aud[24155]=16'hcfa;
aud[24156]=16'hd0f;
aud[24157]=16'hd24;
aud[24158]=16'hd39;
aud[24159]=16'hd4e;
aud[24160]=16'hd63;
aud[24161]=16'hd78;
aud[24162]=16'hd8d;
aud[24163]=16'hda2;
aud[24164]=16'hdb7;
aud[24165]=16'hdcc;
aud[24166]=16'hde1;
aud[24167]=16'hdf6;
aud[24168]=16'he0b;
aud[24169]=16'he20;
aud[24170]=16'he35;
aud[24171]=16'he4a;
aud[24172]=16'he5f;
aud[24173]=16'he74;
aud[24174]=16'he88;
aud[24175]=16'he9d;
aud[24176]=16'heb2;
aud[24177]=16'hec7;
aud[24178]=16'hedc;
aud[24179]=16'hef1;
aud[24180]=16'hf06;
aud[24181]=16'hf1a;
aud[24182]=16'hf2f;
aud[24183]=16'hf44;
aud[24184]=16'hf59;
aud[24185]=16'hf6e;
aud[24186]=16'hf83;
aud[24187]=16'hf97;
aud[24188]=16'hfac;
aud[24189]=16'hfc1;
aud[24190]=16'hfd6;
aud[24191]=16'hfeb;
aud[24192]=16'hfff;
aud[24193]=16'h1014;
aud[24194]=16'h1029;
aud[24195]=16'h103e;
aud[24196]=16'h1052;
aud[24197]=16'h1067;
aud[24198]=16'h107c;
aud[24199]=16'h1090;
aud[24200]=16'h10a5;
aud[24201]=16'h10ba;
aud[24202]=16'h10cf;
aud[24203]=16'h10e3;
aud[24204]=16'h10f8;
aud[24205]=16'h110d;
aud[24206]=16'h1121;
aud[24207]=16'h1136;
aud[24208]=16'h114b;
aud[24209]=16'h115f;
aud[24210]=16'h1174;
aud[24211]=16'h1189;
aud[24212]=16'h119d;
aud[24213]=16'h11b2;
aud[24214]=16'h11c6;
aud[24215]=16'h11db;
aud[24216]=16'h11f0;
aud[24217]=16'h1204;
aud[24218]=16'h1219;
aud[24219]=16'h122d;
aud[24220]=16'h1242;
aud[24221]=16'h1256;
aud[24222]=16'h126b;
aud[24223]=16'h127f;
aud[24224]=16'h1294;
aud[24225]=16'h12a9;
aud[24226]=16'h12bd;
aud[24227]=16'h12d2;
aud[24228]=16'h12e6;
aud[24229]=16'h12fb;
aud[24230]=16'h130f;
aud[24231]=16'h1323;
aud[24232]=16'h1338;
aud[24233]=16'h134c;
aud[24234]=16'h1361;
aud[24235]=16'h1375;
aud[24236]=16'h138a;
aud[24237]=16'h139e;
aud[24238]=16'h13b3;
aud[24239]=16'h13c7;
aud[24240]=16'h13db;
aud[24241]=16'h13f0;
aud[24242]=16'h1404;
aud[24243]=16'h1418;
aud[24244]=16'h142d;
aud[24245]=16'h1441;
aud[24246]=16'h1455;
aud[24247]=16'h146a;
aud[24248]=16'h147e;
aud[24249]=16'h1492;
aud[24250]=16'h14a7;
aud[24251]=16'h14bb;
aud[24252]=16'h14cf;
aud[24253]=16'h14e4;
aud[24254]=16'h14f8;
aud[24255]=16'h150c;
aud[24256]=16'h1520;
aud[24257]=16'h1535;
aud[24258]=16'h1549;
aud[24259]=16'h155d;
aud[24260]=16'h1571;
aud[24261]=16'h1586;
aud[24262]=16'h159a;
aud[24263]=16'h15ae;
aud[24264]=16'h15c2;
aud[24265]=16'h15d6;
aud[24266]=16'h15ea;
aud[24267]=16'h15ff;
aud[24268]=16'h1613;
aud[24269]=16'h1627;
aud[24270]=16'h163b;
aud[24271]=16'h164f;
aud[24272]=16'h1663;
aud[24273]=16'h1677;
aud[24274]=16'h168b;
aud[24275]=16'h169f;
aud[24276]=16'h16b3;
aud[24277]=16'h16c7;
aud[24278]=16'h16db;
aud[24279]=16'h16f0;
aud[24280]=16'h1704;
aud[24281]=16'h1718;
aud[24282]=16'h172c;
aud[24283]=16'h1740;
aud[24284]=16'h1753;
aud[24285]=16'h1767;
aud[24286]=16'h177b;
aud[24287]=16'h178f;
aud[24288]=16'h17a3;
aud[24289]=16'h17b7;
aud[24290]=16'h17cb;
aud[24291]=16'h17df;
aud[24292]=16'h17f3;
aud[24293]=16'h1807;
aud[24294]=16'h181b;
aud[24295]=16'h182f;
aud[24296]=16'h1842;
aud[24297]=16'h1856;
aud[24298]=16'h186a;
aud[24299]=16'h187e;
aud[24300]=16'h1892;
aud[24301]=16'h18a5;
aud[24302]=16'h18b9;
aud[24303]=16'h18cd;
aud[24304]=16'h18e1;
aud[24305]=16'h18f5;
aud[24306]=16'h1908;
aud[24307]=16'h191c;
aud[24308]=16'h1930;
aud[24309]=16'h1943;
aud[24310]=16'h1957;
aud[24311]=16'h196b;
aud[24312]=16'h197f;
aud[24313]=16'h1992;
aud[24314]=16'h19a6;
aud[24315]=16'h19ba;
aud[24316]=16'h19cd;
aud[24317]=16'h19e1;
aud[24318]=16'h19f4;
aud[24319]=16'h1a08;
aud[24320]=16'h1a1c;
aud[24321]=16'h1a2f;
aud[24322]=16'h1a43;
aud[24323]=16'h1a56;
aud[24324]=16'h1a6a;
aud[24325]=16'h1a7d;
aud[24326]=16'h1a91;
aud[24327]=16'h1aa4;
aud[24328]=16'h1ab8;
aud[24329]=16'h1acb;
aud[24330]=16'h1adf;
aud[24331]=16'h1af2;
aud[24332]=16'h1b06;
aud[24333]=16'h1b19;
aud[24334]=16'h1b2d;
aud[24335]=16'h1b40;
aud[24336]=16'h1b53;
aud[24337]=16'h1b67;
aud[24338]=16'h1b7a;
aud[24339]=16'h1b8d;
aud[24340]=16'h1ba1;
aud[24341]=16'h1bb4;
aud[24342]=16'h1bc8;
aud[24343]=16'h1bdb;
aud[24344]=16'h1bee;
aud[24345]=16'h1c01;
aud[24346]=16'h1c15;
aud[24347]=16'h1c28;
aud[24348]=16'h1c3b;
aud[24349]=16'h1c4e;
aud[24350]=16'h1c62;
aud[24351]=16'h1c75;
aud[24352]=16'h1c88;
aud[24353]=16'h1c9b;
aud[24354]=16'h1cae;
aud[24355]=16'h1cc2;
aud[24356]=16'h1cd5;
aud[24357]=16'h1ce8;
aud[24358]=16'h1cfb;
aud[24359]=16'h1d0e;
aud[24360]=16'h1d21;
aud[24361]=16'h1d34;
aud[24362]=16'h1d47;
aud[24363]=16'h1d5b;
aud[24364]=16'h1d6e;
aud[24365]=16'h1d81;
aud[24366]=16'h1d94;
aud[24367]=16'h1da7;
aud[24368]=16'h1dba;
aud[24369]=16'h1dcd;
aud[24370]=16'h1de0;
aud[24371]=16'h1df3;
aud[24372]=16'h1e06;
aud[24373]=16'h1e18;
aud[24374]=16'h1e2b;
aud[24375]=16'h1e3e;
aud[24376]=16'h1e51;
aud[24377]=16'h1e64;
aud[24378]=16'h1e77;
aud[24379]=16'h1e8a;
aud[24380]=16'h1e9d;
aud[24381]=16'h1eaf;
aud[24382]=16'h1ec2;
aud[24383]=16'h1ed5;
aud[24384]=16'h1ee8;
aud[24385]=16'h1efb;
aud[24386]=16'h1f0d;
aud[24387]=16'h1f20;
aud[24388]=16'h1f33;
aud[24389]=16'h1f46;
aud[24390]=16'h1f58;
aud[24391]=16'h1f6b;
aud[24392]=16'h1f7e;
aud[24393]=16'h1f90;
aud[24394]=16'h1fa3;
aud[24395]=16'h1fb6;
aud[24396]=16'h1fc8;
aud[24397]=16'h1fdb;
aud[24398]=16'h1fed;
aud[24399]=16'h2000;
aud[24400]=16'h2013;
aud[24401]=16'h2025;
aud[24402]=16'h2038;
aud[24403]=16'h204a;
aud[24404]=16'h205d;
aud[24405]=16'h206f;
aud[24406]=16'h2082;
aud[24407]=16'h2094;
aud[24408]=16'h20a7;
aud[24409]=16'h20b9;
aud[24410]=16'h20cb;
aud[24411]=16'h20de;
aud[24412]=16'h20f0;
aud[24413]=16'h2103;
aud[24414]=16'h2115;
aud[24415]=16'h2127;
aud[24416]=16'h213a;
aud[24417]=16'h214c;
aud[24418]=16'h215e;
aud[24419]=16'h2171;
aud[24420]=16'h2183;
aud[24421]=16'h2195;
aud[24422]=16'h21a7;
aud[24423]=16'h21ba;
aud[24424]=16'h21cc;
aud[24425]=16'h21de;
aud[24426]=16'h21f0;
aud[24427]=16'h2202;
aud[24428]=16'h2215;
aud[24429]=16'h2227;
aud[24430]=16'h2239;
aud[24431]=16'h224b;
aud[24432]=16'h225d;
aud[24433]=16'h226f;
aud[24434]=16'h2281;
aud[24435]=16'h2293;
aud[24436]=16'h22a5;
aud[24437]=16'h22b7;
aud[24438]=16'h22c9;
aud[24439]=16'h22db;
aud[24440]=16'h22ed;
aud[24441]=16'h22ff;
aud[24442]=16'h2311;
aud[24443]=16'h2323;
aud[24444]=16'h2335;
aud[24445]=16'h2347;
aud[24446]=16'h2359;
aud[24447]=16'h236b;
aud[24448]=16'h237d;
aud[24449]=16'h238e;
aud[24450]=16'h23a0;
aud[24451]=16'h23b2;
aud[24452]=16'h23c4;
aud[24453]=16'h23d6;
aud[24454]=16'h23e7;
aud[24455]=16'h23f9;
aud[24456]=16'h240b;
aud[24457]=16'h241d;
aud[24458]=16'h242e;
aud[24459]=16'h2440;
aud[24460]=16'h2452;
aud[24461]=16'h2463;
aud[24462]=16'h2475;
aud[24463]=16'h2487;
aud[24464]=16'h2498;
aud[24465]=16'h24aa;
aud[24466]=16'h24bb;
aud[24467]=16'h24cd;
aud[24468]=16'h24de;
aud[24469]=16'h24f0;
aud[24470]=16'h2501;
aud[24471]=16'h2513;
aud[24472]=16'h2524;
aud[24473]=16'h2536;
aud[24474]=16'h2547;
aud[24475]=16'h2559;
aud[24476]=16'h256a;
aud[24477]=16'h257c;
aud[24478]=16'h258d;
aud[24479]=16'h259e;
aud[24480]=16'h25b0;
aud[24481]=16'h25c1;
aud[24482]=16'h25d2;
aud[24483]=16'h25e4;
aud[24484]=16'h25f5;
aud[24485]=16'h2606;
aud[24486]=16'h2617;
aud[24487]=16'h2629;
aud[24488]=16'h263a;
aud[24489]=16'h264b;
aud[24490]=16'h265c;
aud[24491]=16'h266d;
aud[24492]=16'h267e;
aud[24493]=16'h2690;
aud[24494]=16'h26a1;
aud[24495]=16'h26b2;
aud[24496]=16'h26c3;
aud[24497]=16'h26d4;
aud[24498]=16'h26e5;
aud[24499]=16'h26f6;
aud[24500]=16'h2707;
aud[24501]=16'h2718;
aud[24502]=16'h2729;
aud[24503]=16'h273a;
aud[24504]=16'h274b;
aud[24505]=16'h275c;
aud[24506]=16'h276d;
aud[24507]=16'h277e;
aud[24508]=16'h278e;
aud[24509]=16'h279f;
aud[24510]=16'h27b0;
aud[24511]=16'h27c1;
aud[24512]=16'h27d2;
aud[24513]=16'h27e2;
aud[24514]=16'h27f3;
aud[24515]=16'h2804;
aud[24516]=16'h2815;
aud[24517]=16'h2825;
aud[24518]=16'h2836;
aud[24519]=16'h2847;
aud[24520]=16'h2857;
aud[24521]=16'h2868;
aud[24522]=16'h2879;
aud[24523]=16'h2889;
aud[24524]=16'h289a;
aud[24525]=16'h28aa;
aud[24526]=16'h28bb;
aud[24527]=16'h28cc;
aud[24528]=16'h28dc;
aud[24529]=16'h28ed;
aud[24530]=16'h28fd;
aud[24531]=16'h290e;
aud[24532]=16'h291e;
aud[24533]=16'h292e;
aud[24534]=16'h293f;
aud[24535]=16'h294f;
aud[24536]=16'h2960;
aud[24537]=16'h2970;
aud[24538]=16'h2980;
aud[24539]=16'h2991;
aud[24540]=16'h29a1;
aud[24541]=16'h29b1;
aud[24542]=16'h29c1;
aud[24543]=16'h29d2;
aud[24544]=16'h29e2;
aud[24545]=16'h29f2;
aud[24546]=16'h2a02;
aud[24547]=16'h2a12;
aud[24548]=16'h2a23;
aud[24549]=16'h2a33;
aud[24550]=16'h2a43;
aud[24551]=16'h2a53;
aud[24552]=16'h2a63;
aud[24553]=16'h2a73;
aud[24554]=16'h2a83;
aud[24555]=16'h2a93;
aud[24556]=16'h2aa3;
aud[24557]=16'h2ab3;
aud[24558]=16'h2ac3;
aud[24559]=16'h2ad3;
aud[24560]=16'h2ae3;
aud[24561]=16'h2af3;
aud[24562]=16'h2b03;
aud[24563]=16'h2b13;
aud[24564]=16'h2b22;
aud[24565]=16'h2b32;
aud[24566]=16'h2b42;
aud[24567]=16'h2b52;
aud[24568]=16'h2b62;
aud[24569]=16'h2b71;
aud[24570]=16'h2b81;
aud[24571]=16'h2b91;
aud[24572]=16'h2ba1;
aud[24573]=16'h2bb0;
aud[24574]=16'h2bc0;
aud[24575]=16'h2bd0;
aud[24576]=16'h2bdf;
aud[24577]=16'h2bef;
aud[24578]=16'h2bfe;
aud[24579]=16'h2c0e;
aud[24580]=16'h2c1e;
aud[24581]=16'h2c2d;
aud[24582]=16'h2c3d;
aud[24583]=16'h2c4c;
aud[24584]=16'h2c5c;
aud[24585]=16'h2c6b;
aud[24586]=16'h2c7a;
aud[24587]=16'h2c8a;
aud[24588]=16'h2c99;
aud[24589]=16'h2ca9;
aud[24590]=16'h2cb8;
aud[24591]=16'h2cc7;
aud[24592]=16'h2cd7;
aud[24593]=16'h2ce6;
aud[24594]=16'h2cf5;
aud[24595]=16'h2d04;
aud[24596]=16'h2d14;
aud[24597]=16'h2d23;
aud[24598]=16'h2d32;
aud[24599]=16'h2d41;
aud[24600]=16'h2d50;
aud[24601]=16'h2d60;
aud[24602]=16'h2d6f;
aud[24603]=16'h2d7e;
aud[24604]=16'h2d8d;
aud[24605]=16'h2d9c;
aud[24606]=16'h2dab;
aud[24607]=16'h2dba;
aud[24608]=16'h2dc9;
aud[24609]=16'h2dd8;
aud[24610]=16'h2de7;
aud[24611]=16'h2df6;
aud[24612]=16'h2e05;
aud[24613]=16'h2e14;
aud[24614]=16'h2e22;
aud[24615]=16'h2e31;
aud[24616]=16'h2e40;
aud[24617]=16'h2e4f;
aud[24618]=16'h2e5e;
aud[24619]=16'h2e6d;
aud[24620]=16'h2e7b;
aud[24621]=16'h2e8a;
aud[24622]=16'h2e99;
aud[24623]=16'h2ea7;
aud[24624]=16'h2eb6;
aud[24625]=16'h2ec5;
aud[24626]=16'h2ed3;
aud[24627]=16'h2ee2;
aud[24628]=16'h2ef1;
aud[24629]=16'h2eff;
aud[24630]=16'h2f0e;
aud[24631]=16'h2f1c;
aud[24632]=16'h2f2b;
aud[24633]=16'h2f39;
aud[24634]=16'h2f48;
aud[24635]=16'h2f56;
aud[24636]=16'h2f65;
aud[24637]=16'h2f73;
aud[24638]=16'h2f81;
aud[24639]=16'h2f90;
aud[24640]=16'h2f9e;
aud[24641]=16'h2fac;
aud[24642]=16'h2fbb;
aud[24643]=16'h2fc9;
aud[24644]=16'h2fd7;
aud[24645]=16'h2fe5;
aud[24646]=16'h2ff4;
aud[24647]=16'h3002;
aud[24648]=16'h3010;
aud[24649]=16'h301e;
aud[24650]=16'h302c;
aud[24651]=16'h303a;
aud[24652]=16'h3048;
aud[24653]=16'h3057;
aud[24654]=16'h3065;
aud[24655]=16'h3073;
aud[24656]=16'h3081;
aud[24657]=16'h308f;
aud[24658]=16'h309d;
aud[24659]=16'h30aa;
aud[24660]=16'h30b8;
aud[24661]=16'h30c6;
aud[24662]=16'h30d4;
aud[24663]=16'h30e2;
aud[24664]=16'h30f0;
aud[24665]=16'h30fe;
aud[24666]=16'h310b;
aud[24667]=16'h3119;
aud[24668]=16'h3127;
aud[24669]=16'h3135;
aud[24670]=16'h3142;
aud[24671]=16'h3150;
aud[24672]=16'h315e;
aud[24673]=16'h316b;
aud[24674]=16'h3179;
aud[24675]=16'h3187;
aud[24676]=16'h3194;
aud[24677]=16'h31a2;
aud[24678]=16'h31af;
aud[24679]=16'h31bd;
aud[24680]=16'h31ca;
aud[24681]=16'h31d8;
aud[24682]=16'h31e5;
aud[24683]=16'h31f3;
aud[24684]=16'h3200;
aud[24685]=16'h320d;
aud[24686]=16'h321b;
aud[24687]=16'h3228;
aud[24688]=16'h3235;
aud[24689]=16'h3243;
aud[24690]=16'h3250;
aud[24691]=16'h325d;
aud[24692]=16'h326a;
aud[24693]=16'h3278;
aud[24694]=16'h3285;
aud[24695]=16'h3292;
aud[24696]=16'h329f;
aud[24697]=16'h32ac;
aud[24698]=16'h32b9;
aud[24699]=16'h32c6;
aud[24700]=16'h32d3;
aud[24701]=16'h32e0;
aud[24702]=16'h32ed;
aud[24703]=16'h32fa;
aud[24704]=16'h3307;
aud[24705]=16'h3314;
aud[24706]=16'h3321;
aud[24707]=16'h332e;
aud[24708]=16'h333b;
aud[24709]=16'h3348;
aud[24710]=16'h3355;
aud[24711]=16'h3361;
aud[24712]=16'h336e;
aud[24713]=16'h337b;
aud[24714]=16'h3388;
aud[24715]=16'h3394;
aud[24716]=16'h33a1;
aud[24717]=16'h33ae;
aud[24718]=16'h33ba;
aud[24719]=16'h33c7;
aud[24720]=16'h33d4;
aud[24721]=16'h33e0;
aud[24722]=16'h33ed;
aud[24723]=16'h33f9;
aud[24724]=16'h3406;
aud[24725]=16'h3412;
aud[24726]=16'h341f;
aud[24727]=16'h342b;
aud[24728]=16'h3437;
aud[24729]=16'h3444;
aud[24730]=16'h3450;
aud[24731]=16'h345d;
aud[24732]=16'h3469;
aud[24733]=16'h3475;
aud[24734]=16'h3481;
aud[24735]=16'h348e;
aud[24736]=16'h349a;
aud[24737]=16'h34a6;
aud[24738]=16'h34b2;
aud[24739]=16'h34be;
aud[24740]=16'h34cb;
aud[24741]=16'h34d7;
aud[24742]=16'h34e3;
aud[24743]=16'h34ef;
aud[24744]=16'h34fb;
aud[24745]=16'h3507;
aud[24746]=16'h3513;
aud[24747]=16'h351f;
aud[24748]=16'h352b;
aud[24749]=16'h3537;
aud[24750]=16'h3543;
aud[24751]=16'h354f;
aud[24752]=16'h355a;
aud[24753]=16'h3566;
aud[24754]=16'h3572;
aud[24755]=16'h357e;
aud[24756]=16'h358a;
aud[24757]=16'h3595;
aud[24758]=16'h35a1;
aud[24759]=16'h35ad;
aud[24760]=16'h35b8;
aud[24761]=16'h35c4;
aud[24762]=16'h35d0;
aud[24763]=16'h35db;
aud[24764]=16'h35e7;
aud[24765]=16'h35f2;
aud[24766]=16'h35fe;
aud[24767]=16'h3609;
aud[24768]=16'h3615;
aud[24769]=16'h3620;
aud[24770]=16'h362c;
aud[24771]=16'h3637;
aud[24772]=16'h3643;
aud[24773]=16'h364e;
aud[24774]=16'h3659;
aud[24775]=16'h3665;
aud[24776]=16'h3670;
aud[24777]=16'h367b;
aud[24778]=16'h3686;
aud[24779]=16'h3692;
aud[24780]=16'h369d;
aud[24781]=16'h36a8;
aud[24782]=16'h36b3;
aud[24783]=16'h36be;
aud[24784]=16'h36c9;
aud[24785]=16'h36d4;
aud[24786]=16'h36e0;
aud[24787]=16'h36eb;
aud[24788]=16'h36f6;
aud[24789]=16'h3701;
aud[24790]=16'h370b;
aud[24791]=16'h3716;
aud[24792]=16'h3721;
aud[24793]=16'h372c;
aud[24794]=16'h3737;
aud[24795]=16'h3742;
aud[24796]=16'h374d;
aud[24797]=16'h3757;
aud[24798]=16'h3762;
aud[24799]=16'h376d;
aud[24800]=16'h3778;
aud[24801]=16'h3782;
aud[24802]=16'h378d;
aud[24803]=16'h3798;
aud[24804]=16'h37a2;
aud[24805]=16'h37ad;
aud[24806]=16'h37b7;
aud[24807]=16'h37c2;
aud[24808]=16'h37cc;
aud[24809]=16'h37d7;
aud[24810]=16'h37e1;
aud[24811]=16'h37ec;
aud[24812]=16'h37f6;
aud[24813]=16'h3801;
aud[24814]=16'h380b;
aud[24815]=16'h3815;
aud[24816]=16'h3820;
aud[24817]=16'h382a;
aud[24818]=16'h3834;
aud[24819]=16'h383f;
aud[24820]=16'h3849;
aud[24821]=16'h3853;
aud[24822]=16'h385d;
aud[24823]=16'h3867;
aud[24824]=16'h3871;
aud[24825]=16'h387b;
aud[24826]=16'h3886;
aud[24827]=16'h3890;
aud[24828]=16'h389a;
aud[24829]=16'h38a4;
aud[24830]=16'h38ae;
aud[24831]=16'h38b8;
aud[24832]=16'h38c1;
aud[24833]=16'h38cb;
aud[24834]=16'h38d5;
aud[24835]=16'h38df;
aud[24836]=16'h38e9;
aud[24837]=16'h38f3;
aud[24838]=16'h38fd;
aud[24839]=16'h3906;
aud[24840]=16'h3910;
aud[24841]=16'h391a;
aud[24842]=16'h3923;
aud[24843]=16'h392d;
aud[24844]=16'h3937;
aud[24845]=16'h3940;
aud[24846]=16'h394a;
aud[24847]=16'h3953;
aud[24848]=16'h395d;
aud[24849]=16'h3966;
aud[24850]=16'h3970;
aud[24851]=16'h3979;
aud[24852]=16'h3983;
aud[24853]=16'h398c;
aud[24854]=16'h3995;
aud[24855]=16'h399f;
aud[24856]=16'h39a8;
aud[24857]=16'h39b1;
aud[24858]=16'h39bb;
aud[24859]=16'h39c4;
aud[24860]=16'h39cd;
aud[24861]=16'h39d6;
aud[24862]=16'h39e0;
aud[24863]=16'h39e9;
aud[24864]=16'h39f2;
aud[24865]=16'h39fb;
aud[24866]=16'h3a04;
aud[24867]=16'h3a0d;
aud[24868]=16'h3a16;
aud[24869]=16'h3a1f;
aud[24870]=16'h3a28;
aud[24871]=16'h3a31;
aud[24872]=16'h3a3a;
aud[24873]=16'h3a43;
aud[24874]=16'h3a4c;
aud[24875]=16'h3a54;
aud[24876]=16'h3a5d;
aud[24877]=16'h3a66;
aud[24878]=16'h3a6f;
aud[24879]=16'h3a78;
aud[24880]=16'h3a80;
aud[24881]=16'h3a89;
aud[24882]=16'h3a92;
aud[24883]=16'h3a9a;
aud[24884]=16'h3aa3;
aud[24885]=16'h3aab;
aud[24886]=16'h3ab4;
aud[24887]=16'h3abc;
aud[24888]=16'h3ac5;
aud[24889]=16'h3acd;
aud[24890]=16'h3ad6;
aud[24891]=16'h3ade;
aud[24892]=16'h3ae7;
aud[24893]=16'h3aef;
aud[24894]=16'h3af7;
aud[24895]=16'h3b00;
aud[24896]=16'h3b08;
aud[24897]=16'h3b10;
aud[24898]=16'h3b19;
aud[24899]=16'h3b21;
aud[24900]=16'h3b29;
aud[24901]=16'h3b31;
aud[24902]=16'h3b39;
aud[24903]=16'h3b41;
aud[24904]=16'h3b4a;
aud[24905]=16'h3b52;
aud[24906]=16'h3b5a;
aud[24907]=16'h3b62;
aud[24908]=16'h3b6a;
aud[24909]=16'h3b72;
aud[24910]=16'h3b7a;
aud[24911]=16'h3b81;
aud[24912]=16'h3b89;
aud[24913]=16'h3b91;
aud[24914]=16'h3b99;
aud[24915]=16'h3ba1;
aud[24916]=16'h3ba9;
aud[24917]=16'h3bb0;
aud[24918]=16'h3bb8;
aud[24919]=16'h3bc0;
aud[24920]=16'h3bc7;
aud[24921]=16'h3bcf;
aud[24922]=16'h3bd7;
aud[24923]=16'h3bde;
aud[24924]=16'h3be6;
aud[24925]=16'h3bed;
aud[24926]=16'h3bf5;
aud[24927]=16'h3bfc;
aud[24928]=16'h3c04;
aud[24929]=16'h3c0b;
aud[24930]=16'h3c13;
aud[24931]=16'h3c1a;
aud[24932]=16'h3c21;
aud[24933]=16'h3c29;
aud[24934]=16'h3c30;
aud[24935]=16'h3c37;
aud[24936]=16'h3c3f;
aud[24937]=16'h3c46;
aud[24938]=16'h3c4d;
aud[24939]=16'h3c54;
aud[24940]=16'h3c5b;
aud[24941]=16'h3c63;
aud[24942]=16'h3c6a;
aud[24943]=16'h3c71;
aud[24944]=16'h3c78;
aud[24945]=16'h3c7f;
aud[24946]=16'h3c86;
aud[24947]=16'h3c8d;
aud[24948]=16'h3c94;
aud[24949]=16'h3c9b;
aud[24950]=16'h3ca1;
aud[24951]=16'h3ca8;
aud[24952]=16'h3caf;
aud[24953]=16'h3cb6;
aud[24954]=16'h3cbd;
aud[24955]=16'h3cc3;
aud[24956]=16'h3cca;
aud[24957]=16'h3cd1;
aud[24958]=16'h3cd7;
aud[24959]=16'h3cde;
aud[24960]=16'h3ce5;
aud[24961]=16'h3ceb;
aud[24962]=16'h3cf2;
aud[24963]=16'h3cf8;
aud[24964]=16'h3cff;
aud[24965]=16'h3d05;
aud[24966]=16'h3d0c;
aud[24967]=16'h3d12;
aud[24968]=16'h3d19;
aud[24969]=16'h3d1f;
aud[24970]=16'h3d25;
aud[24971]=16'h3d2c;
aud[24972]=16'h3d32;
aud[24973]=16'h3d38;
aud[24974]=16'h3d3f;
aud[24975]=16'h3d45;
aud[24976]=16'h3d4b;
aud[24977]=16'h3d51;
aud[24978]=16'h3d57;
aud[24979]=16'h3d5d;
aud[24980]=16'h3d63;
aud[24981]=16'h3d69;
aud[24982]=16'h3d6f;
aud[24983]=16'h3d75;
aud[24984]=16'h3d7b;
aud[24985]=16'h3d81;
aud[24986]=16'h3d87;
aud[24987]=16'h3d8d;
aud[24988]=16'h3d93;
aud[24989]=16'h3d99;
aud[24990]=16'h3d9f;
aud[24991]=16'h3da4;
aud[24992]=16'h3daa;
aud[24993]=16'h3db0;
aud[24994]=16'h3db6;
aud[24995]=16'h3dbb;
aud[24996]=16'h3dc1;
aud[24997]=16'h3dc7;
aud[24998]=16'h3dcc;
aud[24999]=16'h3dd2;
aud[25000]=16'h3dd7;
aud[25001]=16'h3ddd;
aud[25002]=16'h3de2;
aud[25003]=16'h3de8;
aud[25004]=16'h3ded;
aud[25005]=16'h3df3;
aud[25006]=16'h3df8;
aud[25007]=16'h3dfd;
aud[25008]=16'h3e03;
aud[25009]=16'h3e08;
aud[25010]=16'h3e0d;
aud[25011]=16'h3e12;
aud[25012]=16'h3e18;
aud[25013]=16'h3e1d;
aud[25014]=16'h3e22;
aud[25015]=16'h3e27;
aud[25016]=16'h3e2c;
aud[25017]=16'h3e31;
aud[25018]=16'h3e36;
aud[25019]=16'h3e3b;
aud[25020]=16'h3e40;
aud[25021]=16'h3e45;
aud[25022]=16'h3e4a;
aud[25023]=16'h3e4f;
aud[25024]=16'h3e54;
aud[25025]=16'h3e59;
aud[25026]=16'h3e5e;
aud[25027]=16'h3e62;
aud[25028]=16'h3e67;
aud[25029]=16'h3e6c;
aud[25030]=16'h3e71;
aud[25031]=16'h3e75;
aud[25032]=16'h3e7a;
aud[25033]=16'h3e7f;
aud[25034]=16'h3e83;
aud[25035]=16'h3e88;
aud[25036]=16'h3e8c;
aud[25037]=16'h3e91;
aud[25038]=16'h3e95;
aud[25039]=16'h3e9a;
aud[25040]=16'h3e9e;
aud[25041]=16'h3ea3;
aud[25042]=16'h3ea7;
aud[25043]=16'h3eac;
aud[25044]=16'h3eb0;
aud[25045]=16'h3eb4;
aud[25046]=16'h3eb9;
aud[25047]=16'h3ebd;
aud[25048]=16'h3ec1;
aud[25049]=16'h3ec5;
aud[25050]=16'h3ec9;
aud[25051]=16'h3ecd;
aud[25052]=16'h3ed2;
aud[25053]=16'h3ed6;
aud[25054]=16'h3eda;
aud[25055]=16'h3ede;
aud[25056]=16'h3ee2;
aud[25057]=16'h3ee6;
aud[25058]=16'h3eea;
aud[25059]=16'h3eee;
aud[25060]=16'h3ef2;
aud[25061]=16'h3ef5;
aud[25062]=16'h3ef9;
aud[25063]=16'h3efd;
aud[25064]=16'h3f01;
aud[25065]=16'h3f05;
aud[25066]=16'h3f08;
aud[25067]=16'h3f0c;
aud[25068]=16'h3f10;
aud[25069]=16'h3f13;
aud[25070]=16'h3f17;
aud[25071]=16'h3f1b;
aud[25072]=16'h3f1e;
aud[25073]=16'h3f22;
aud[25074]=16'h3f25;
aud[25075]=16'h3f29;
aud[25076]=16'h3f2c;
aud[25077]=16'h3f30;
aud[25078]=16'h3f33;
aud[25079]=16'h3f36;
aud[25080]=16'h3f3a;
aud[25081]=16'h3f3d;
aud[25082]=16'h3f40;
aud[25083]=16'h3f43;
aud[25084]=16'h3f47;
aud[25085]=16'h3f4a;
aud[25086]=16'h3f4d;
aud[25087]=16'h3f50;
aud[25088]=16'h3f53;
aud[25089]=16'h3f56;
aud[25090]=16'h3f5a;
aud[25091]=16'h3f5d;
aud[25092]=16'h3f60;
aud[25093]=16'h3f63;
aud[25094]=16'h3f65;
aud[25095]=16'h3f68;
aud[25096]=16'h3f6b;
aud[25097]=16'h3f6e;
aud[25098]=16'h3f71;
aud[25099]=16'h3f74;
aud[25100]=16'h3f77;
aud[25101]=16'h3f79;
aud[25102]=16'h3f7c;
aud[25103]=16'h3f7f;
aud[25104]=16'h3f81;
aud[25105]=16'h3f84;
aud[25106]=16'h3f87;
aud[25107]=16'h3f89;
aud[25108]=16'h3f8c;
aud[25109]=16'h3f8e;
aud[25110]=16'h3f91;
aud[25111]=16'h3f93;
aud[25112]=16'h3f96;
aud[25113]=16'h3f98;
aud[25114]=16'h3f9b;
aud[25115]=16'h3f9d;
aud[25116]=16'h3f9f;
aud[25117]=16'h3fa2;
aud[25118]=16'h3fa4;
aud[25119]=16'h3fa6;
aud[25120]=16'h3fa8;
aud[25121]=16'h3fab;
aud[25122]=16'h3fad;
aud[25123]=16'h3faf;
aud[25124]=16'h3fb1;
aud[25125]=16'h3fb3;
aud[25126]=16'h3fb5;
aud[25127]=16'h3fb7;
aud[25128]=16'h3fb9;
aud[25129]=16'h3fbb;
aud[25130]=16'h3fbd;
aud[25131]=16'h3fbf;
aud[25132]=16'h3fc1;
aud[25133]=16'h3fc3;
aud[25134]=16'h3fc5;
aud[25135]=16'h3fc7;
aud[25136]=16'h3fc8;
aud[25137]=16'h3fca;
aud[25138]=16'h3fcc;
aud[25139]=16'h3fcd;
aud[25140]=16'h3fcf;
aud[25141]=16'h3fd1;
aud[25142]=16'h3fd2;
aud[25143]=16'h3fd4;
aud[25144]=16'h3fd6;
aud[25145]=16'h3fd7;
aud[25146]=16'h3fd9;
aud[25147]=16'h3fda;
aud[25148]=16'h3fdc;
aud[25149]=16'h3fdd;
aud[25150]=16'h3fde;
aud[25151]=16'h3fe0;
aud[25152]=16'h3fe1;
aud[25153]=16'h3fe2;
aud[25154]=16'h3fe4;
aud[25155]=16'h3fe5;
aud[25156]=16'h3fe6;
aud[25157]=16'h3fe7;
aud[25158]=16'h3fe8;
aud[25159]=16'h3fea;
aud[25160]=16'h3feb;
aud[25161]=16'h3fec;
aud[25162]=16'h3fed;
aud[25163]=16'h3fee;
aud[25164]=16'h3fef;
aud[25165]=16'h3ff0;
aud[25166]=16'h3ff1;
aud[25167]=16'h3ff2;
aud[25168]=16'h3ff3;
aud[25169]=16'h3ff3;
aud[25170]=16'h3ff4;
aud[25171]=16'h3ff5;
aud[25172]=16'h3ff6;
aud[25173]=16'h3ff7;
aud[25174]=16'h3ff7;
aud[25175]=16'h3ff8;
aud[25176]=16'h3ff9;
aud[25177]=16'h3ff9;
aud[25178]=16'h3ffa;
aud[25179]=16'h3ffa;
aud[25180]=16'h3ffb;
aud[25181]=16'h3ffb;
aud[25182]=16'h3ffc;
aud[25183]=16'h3ffc;
aud[25184]=16'h3ffd;
aud[25185]=16'h3ffd;
aud[25186]=16'h3ffe;
aud[25187]=16'h3ffe;
aud[25188]=16'h3ffe;
aud[25189]=16'h3fff;
aud[25190]=16'h3fff;
aud[25191]=16'h3fff;
aud[25192]=16'h3fff;
aud[25193]=16'h3fff;
aud[25194]=16'h4000;
aud[25195]=16'h4000;
aud[25196]=16'h4000;
aud[25197]=16'h4000;
aud[25198]=16'h4000;
aud[25199]=16'h4000;
aud[25200]=16'h4000;
aud[25201]=16'h4000;
aud[25202]=16'h4000;
aud[25203]=16'h4000;
aud[25204]=16'h4000;
aud[25205]=16'h3fff;
aud[25206]=16'h3fff;
aud[25207]=16'h3fff;
aud[25208]=16'h3fff;
aud[25209]=16'h3fff;
aud[25210]=16'h3ffe;
aud[25211]=16'h3ffe;
aud[25212]=16'h3ffe;
aud[25213]=16'h3ffd;
aud[25214]=16'h3ffd;
aud[25215]=16'h3ffc;
aud[25216]=16'h3ffc;
aud[25217]=16'h3ffb;
aud[25218]=16'h3ffb;
aud[25219]=16'h3ffa;
aud[25220]=16'h3ffa;
aud[25221]=16'h3ff9;
aud[25222]=16'h3ff9;
aud[25223]=16'h3ff8;
aud[25224]=16'h3ff7;
aud[25225]=16'h3ff7;
aud[25226]=16'h3ff6;
aud[25227]=16'h3ff5;
aud[25228]=16'h3ff4;
aud[25229]=16'h3ff3;
aud[25230]=16'h3ff3;
aud[25231]=16'h3ff2;
aud[25232]=16'h3ff1;
aud[25233]=16'h3ff0;
aud[25234]=16'h3fef;
aud[25235]=16'h3fee;
aud[25236]=16'h3fed;
aud[25237]=16'h3fec;
aud[25238]=16'h3feb;
aud[25239]=16'h3fea;
aud[25240]=16'h3fe8;
aud[25241]=16'h3fe7;
aud[25242]=16'h3fe6;
aud[25243]=16'h3fe5;
aud[25244]=16'h3fe4;
aud[25245]=16'h3fe2;
aud[25246]=16'h3fe1;
aud[25247]=16'h3fe0;
aud[25248]=16'h3fde;
aud[25249]=16'h3fdd;
aud[25250]=16'h3fdc;
aud[25251]=16'h3fda;
aud[25252]=16'h3fd9;
aud[25253]=16'h3fd7;
aud[25254]=16'h3fd6;
aud[25255]=16'h3fd4;
aud[25256]=16'h3fd2;
aud[25257]=16'h3fd1;
aud[25258]=16'h3fcf;
aud[25259]=16'h3fcd;
aud[25260]=16'h3fcc;
aud[25261]=16'h3fca;
aud[25262]=16'h3fc8;
aud[25263]=16'h3fc7;
aud[25264]=16'h3fc5;
aud[25265]=16'h3fc3;
aud[25266]=16'h3fc1;
aud[25267]=16'h3fbf;
aud[25268]=16'h3fbd;
aud[25269]=16'h3fbb;
aud[25270]=16'h3fb9;
aud[25271]=16'h3fb7;
aud[25272]=16'h3fb5;
aud[25273]=16'h3fb3;
aud[25274]=16'h3fb1;
aud[25275]=16'h3faf;
aud[25276]=16'h3fad;
aud[25277]=16'h3fab;
aud[25278]=16'h3fa8;
aud[25279]=16'h3fa6;
aud[25280]=16'h3fa4;
aud[25281]=16'h3fa2;
aud[25282]=16'h3f9f;
aud[25283]=16'h3f9d;
aud[25284]=16'h3f9b;
aud[25285]=16'h3f98;
aud[25286]=16'h3f96;
aud[25287]=16'h3f93;
aud[25288]=16'h3f91;
aud[25289]=16'h3f8e;
aud[25290]=16'h3f8c;
aud[25291]=16'h3f89;
aud[25292]=16'h3f87;
aud[25293]=16'h3f84;
aud[25294]=16'h3f81;
aud[25295]=16'h3f7f;
aud[25296]=16'h3f7c;
aud[25297]=16'h3f79;
aud[25298]=16'h3f77;
aud[25299]=16'h3f74;
aud[25300]=16'h3f71;
aud[25301]=16'h3f6e;
aud[25302]=16'h3f6b;
aud[25303]=16'h3f68;
aud[25304]=16'h3f65;
aud[25305]=16'h3f63;
aud[25306]=16'h3f60;
aud[25307]=16'h3f5d;
aud[25308]=16'h3f5a;
aud[25309]=16'h3f56;
aud[25310]=16'h3f53;
aud[25311]=16'h3f50;
aud[25312]=16'h3f4d;
aud[25313]=16'h3f4a;
aud[25314]=16'h3f47;
aud[25315]=16'h3f43;
aud[25316]=16'h3f40;
aud[25317]=16'h3f3d;
aud[25318]=16'h3f3a;
aud[25319]=16'h3f36;
aud[25320]=16'h3f33;
aud[25321]=16'h3f30;
aud[25322]=16'h3f2c;
aud[25323]=16'h3f29;
aud[25324]=16'h3f25;
aud[25325]=16'h3f22;
aud[25326]=16'h3f1e;
aud[25327]=16'h3f1b;
aud[25328]=16'h3f17;
aud[25329]=16'h3f13;
aud[25330]=16'h3f10;
aud[25331]=16'h3f0c;
aud[25332]=16'h3f08;
aud[25333]=16'h3f05;
aud[25334]=16'h3f01;
aud[25335]=16'h3efd;
aud[25336]=16'h3ef9;
aud[25337]=16'h3ef5;
aud[25338]=16'h3ef2;
aud[25339]=16'h3eee;
aud[25340]=16'h3eea;
aud[25341]=16'h3ee6;
aud[25342]=16'h3ee2;
aud[25343]=16'h3ede;
aud[25344]=16'h3eda;
aud[25345]=16'h3ed6;
aud[25346]=16'h3ed2;
aud[25347]=16'h3ecd;
aud[25348]=16'h3ec9;
aud[25349]=16'h3ec5;
aud[25350]=16'h3ec1;
aud[25351]=16'h3ebd;
aud[25352]=16'h3eb9;
aud[25353]=16'h3eb4;
aud[25354]=16'h3eb0;
aud[25355]=16'h3eac;
aud[25356]=16'h3ea7;
aud[25357]=16'h3ea3;
aud[25358]=16'h3e9e;
aud[25359]=16'h3e9a;
aud[25360]=16'h3e95;
aud[25361]=16'h3e91;
aud[25362]=16'h3e8c;
aud[25363]=16'h3e88;
aud[25364]=16'h3e83;
aud[25365]=16'h3e7f;
aud[25366]=16'h3e7a;
aud[25367]=16'h3e75;
aud[25368]=16'h3e71;
aud[25369]=16'h3e6c;
aud[25370]=16'h3e67;
aud[25371]=16'h3e62;
aud[25372]=16'h3e5e;
aud[25373]=16'h3e59;
aud[25374]=16'h3e54;
aud[25375]=16'h3e4f;
aud[25376]=16'h3e4a;
aud[25377]=16'h3e45;
aud[25378]=16'h3e40;
aud[25379]=16'h3e3b;
aud[25380]=16'h3e36;
aud[25381]=16'h3e31;
aud[25382]=16'h3e2c;
aud[25383]=16'h3e27;
aud[25384]=16'h3e22;
aud[25385]=16'h3e1d;
aud[25386]=16'h3e18;
aud[25387]=16'h3e12;
aud[25388]=16'h3e0d;
aud[25389]=16'h3e08;
aud[25390]=16'h3e03;
aud[25391]=16'h3dfd;
aud[25392]=16'h3df8;
aud[25393]=16'h3df3;
aud[25394]=16'h3ded;
aud[25395]=16'h3de8;
aud[25396]=16'h3de2;
aud[25397]=16'h3ddd;
aud[25398]=16'h3dd7;
aud[25399]=16'h3dd2;
aud[25400]=16'h3dcc;
aud[25401]=16'h3dc7;
aud[25402]=16'h3dc1;
aud[25403]=16'h3dbb;
aud[25404]=16'h3db6;
aud[25405]=16'h3db0;
aud[25406]=16'h3daa;
aud[25407]=16'h3da4;
aud[25408]=16'h3d9f;
aud[25409]=16'h3d99;
aud[25410]=16'h3d93;
aud[25411]=16'h3d8d;
aud[25412]=16'h3d87;
aud[25413]=16'h3d81;
aud[25414]=16'h3d7b;
aud[25415]=16'h3d75;
aud[25416]=16'h3d6f;
aud[25417]=16'h3d69;
aud[25418]=16'h3d63;
aud[25419]=16'h3d5d;
aud[25420]=16'h3d57;
aud[25421]=16'h3d51;
aud[25422]=16'h3d4b;
aud[25423]=16'h3d45;
aud[25424]=16'h3d3f;
aud[25425]=16'h3d38;
aud[25426]=16'h3d32;
aud[25427]=16'h3d2c;
aud[25428]=16'h3d25;
aud[25429]=16'h3d1f;
aud[25430]=16'h3d19;
aud[25431]=16'h3d12;
aud[25432]=16'h3d0c;
aud[25433]=16'h3d05;
aud[25434]=16'h3cff;
aud[25435]=16'h3cf8;
aud[25436]=16'h3cf2;
aud[25437]=16'h3ceb;
aud[25438]=16'h3ce5;
aud[25439]=16'h3cde;
aud[25440]=16'h3cd7;
aud[25441]=16'h3cd1;
aud[25442]=16'h3cca;
aud[25443]=16'h3cc3;
aud[25444]=16'h3cbd;
aud[25445]=16'h3cb6;
aud[25446]=16'h3caf;
aud[25447]=16'h3ca8;
aud[25448]=16'h3ca1;
aud[25449]=16'h3c9b;
aud[25450]=16'h3c94;
aud[25451]=16'h3c8d;
aud[25452]=16'h3c86;
aud[25453]=16'h3c7f;
aud[25454]=16'h3c78;
aud[25455]=16'h3c71;
aud[25456]=16'h3c6a;
aud[25457]=16'h3c63;
aud[25458]=16'h3c5b;
aud[25459]=16'h3c54;
aud[25460]=16'h3c4d;
aud[25461]=16'h3c46;
aud[25462]=16'h3c3f;
aud[25463]=16'h3c37;
aud[25464]=16'h3c30;
aud[25465]=16'h3c29;
aud[25466]=16'h3c21;
aud[25467]=16'h3c1a;
aud[25468]=16'h3c13;
aud[25469]=16'h3c0b;
aud[25470]=16'h3c04;
aud[25471]=16'h3bfc;
aud[25472]=16'h3bf5;
aud[25473]=16'h3bed;
aud[25474]=16'h3be6;
aud[25475]=16'h3bde;
aud[25476]=16'h3bd7;
aud[25477]=16'h3bcf;
aud[25478]=16'h3bc7;
aud[25479]=16'h3bc0;
aud[25480]=16'h3bb8;
aud[25481]=16'h3bb0;
aud[25482]=16'h3ba9;
aud[25483]=16'h3ba1;
aud[25484]=16'h3b99;
aud[25485]=16'h3b91;
aud[25486]=16'h3b89;
aud[25487]=16'h3b81;
aud[25488]=16'h3b7a;
aud[25489]=16'h3b72;
aud[25490]=16'h3b6a;
aud[25491]=16'h3b62;
aud[25492]=16'h3b5a;
aud[25493]=16'h3b52;
aud[25494]=16'h3b4a;
aud[25495]=16'h3b41;
aud[25496]=16'h3b39;
aud[25497]=16'h3b31;
aud[25498]=16'h3b29;
aud[25499]=16'h3b21;
aud[25500]=16'h3b19;
aud[25501]=16'h3b10;
aud[25502]=16'h3b08;
aud[25503]=16'h3b00;
aud[25504]=16'h3af7;
aud[25505]=16'h3aef;
aud[25506]=16'h3ae7;
aud[25507]=16'h3ade;
aud[25508]=16'h3ad6;
aud[25509]=16'h3acd;
aud[25510]=16'h3ac5;
aud[25511]=16'h3abc;
aud[25512]=16'h3ab4;
aud[25513]=16'h3aab;
aud[25514]=16'h3aa3;
aud[25515]=16'h3a9a;
aud[25516]=16'h3a92;
aud[25517]=16'h3a89;
aud[25518]=16'h3a80;
aud[25519]=16'h3a78;
aud[25520]=16'h3a6f;
aud[25521]=16'h3a66;
aud[25522]=16'h3a5d;
aud[25523]=16'h3a54;
aud[25524]=16'h3a4c;
aud[25525]=16'h3a43;
aud[25526]=16'h3a3a;
aud[25527]=16'h3a31;
aud[25528]=16'h3a28;
aud[25529]=16'h3a1f;
aud[25530]=16'h3a16;
aud[25531]=16'h3a0d;
aud[25532]=16'h3a04;
aud[25533]=16'h39fb;
aud[25534]=16'h39f2;
aud[25535]=16'h39e9;
aud[25536]=16'h39e0;
aud[25537]=16'h39d6;
aud[25538]=16'h39cd;
aud[25539]=16'h39c4;
aud[25540]=16'h39bb;
aud[25541]=16'h39b1;
aud[25542]=16'h39a8;
aud[25543]=16'h399f;
aud[25544]=16'h3995;
aud[25545]=16'h398c;
aud[25546]=16'h3983;
aud[25547]=16'h3979;
aud[25548]=16'h3970;
aud[25549]=16'h3966;
aud[25550]=16'h395d;
aud[25551]=16'h3953;
aud[25552]=16'h394a;
aud[25553]=16'h3940;
aud[25554]=16'h3937;
aud[25555]=16'h392d;
aud[25556]=16'h3923;
aud[25557]=16'h391a;
aud[25558]=16'h3910;
aud[25559]=16'h3906;
aud[25560]=16'h38fd;
aud[25561]=16'h38f3;
aud[25562]=16'h38e9;
aud[25563]=16'h38df;
aud[25564]=16'h38d5;
aud[25565]=16'h38cb;
aud[25566]=16'h38c1;
aud[25567]=16'h38b8;
aud[25568]=16'h38ae;
aud[25569]=16'h38a4;
aud[25570]=16'h389a;
aud[25571]=16'h3890;
aud[25572]=16'h3886;
aud[25573]=16'h387b;
aud[25574]=16'h3871;
aud[25575]=16'h3867;
aud[25576]=16'h385d;
aud[25577]=16'h3853;
aud[25578]=16'h3849;
aud[25579]=16'h383f;
aud[25580]=16'h3834;
aud[25581]=16'h382a;
aud[25582]=16'h3820;
aud[25583]=16'h3815;
aud[25584]=16'h380b;
aud[25585]=16'h3801;
aud[25586]=16'h37f6;
aud[25587]=16'h37ec;
aud[25588]=16'h37e1;
aud[25589]=16'h37d7;
aud[25590]=16'h37cc;
aud[25591]=16'h37c2;
aud[25592]=16'h37b7;
aud[25593]=16'h37ad;
aud[25594]=16'h37a2;
aud[25595]=16'h3798;
aud[25596]=16'h378d;
aud[25597]=16'h3782;
aud[25598]=16'h3778;
aud[25599]=16'h376d;
aud[25600]=16'h3762;
aud[25601]=16'h3757;
aud[25602]=16'h374d;
aud[25603]=16'h3742;
aud[25604]=16'h3737;
aud[25605]=16'h372c;
aud[25606]=16'h3721;
aud[25607]=16'h3716;
aud[25608]=16'h370b;
aud[25609]=16'h3701;
aud[25610]=16'h36f6;
aud[25611]=16'h36eb;
aud[25612]=16'h36e0;
aud[25613]=16'h36d4;
aud[25614]=16'h36c9;
aud[25615]=16'h36be;
aud[25616]=16'h36b3;
aud[25617]=16'h36a8;
aud[25618]=16'h369d;
aud[25619]=16'h3692;
aud[25620]=16'h3686;
aud[25621]=16'h367b;
aud[25622]=16'h3670;
aud[25623]=16'h3665;
aud[25624]=16'h3659;
aud[25625]=16'h364e;
aud[25626]=16'h3643;
aud[25627]=16'h3637;
aud[25628]=16'h362c;
aud[25629]=16'h3620;
aud[25630]=16'h3615;
aud[25631]=16'h3609;
aud[25632]=16'h35fe;
aud[25633]=16'h35f2;
aud[25634]=16'h35e7;
aud[25635]=16'h35db;
aud[25636]=16'h35d0;
aud[25637]=16'h35c4;
aud[25638]=16'h35b8;
aud[25639]=16'h35ad;
aud[25640]=16'h35a1;
aud[25641]=16'h3595;
aud[25642]=16'h358a;
aud[25643]=16'h357e;
aud[25644]=16'h3572;
aud[25645]=16'h3566;
aud[25646]=16'h355a;
aud[25647]=16'h354f;
aud[25648]=16'h3543;
aud[25649]=16'h3537;
aud[25650]=16'h352b;
aud[25651]=16'h351f;
aud[25652]=16'h3513;
aud[25653]=16'h3507;
aud[25654]=16'h34fb;
aud[25655]=16'h34ef;
aud[25656]=16'h34e3;
aud[25657]=16'h34d7;
aud[25658]=16'h34cb;
aud[25659]=16'h34be;
aud[25660]=16'h34b2;
aud[25661]=16'h34a6;
aud[25662]=16'h349a;
aud[25663]=16'h348e;
aud[25664]=16'h3481;
aud[25665]=16'h3475;
aud[25666]=16'h3469;
aud[25667]=16'h345d;
aud[25668]=16'h3450;
aud[25669]=16'h3444;
aud[25670]=16'h3437;
aud[25671]=16'h342b;
aud[25672]=16'h341f;
aud[25673]=16'h3412;
aud[25674]=16'h3406;
aud[25675]=16'h33f9;
aud[25676]=16'h33ed;
aud[25677]=16'h33e0;
aud[25678]=16'h33d4;
aud[25679]=16'h33c7;
aud[25680]=16'h33ba;
aud[25681]=16'h33ae;
aud[25682]=16'h33a1;
aud[25683]=16'h3394;
aud[25684]=16'h3388;
aud[25685]=16'h337b;
aud[25686]=16'h336e;
aud[25687]=16'h3361;
aud[25688]=16'h3355;
aud[25689]=16'h3348;
aud[25690]=16'h333b;
aud[25691]=16'h332e;
aud[25692]=16'h3321;
aud[25693]=16'h3314;
aud[25694]=16'h3307;
aud[25695]=16'h32fa;
aud[25696]=16'h32ed;
aud[25697]=16'h32e0;
aud[25698]=16'h32d3;
aud[25699]=16'h32c6;
aud[25700]=16'h32b9;
aud[25701]=16'h32ac;
aud[25702]=16'h329f;
aud[25703]=16'h3292;
aud[25704]=16'h3285;
aud[25705]=16'h3278;
aud[25706]=16'h326a;
aud[25707]=16'h325d;
aud[25708]=16'h3250;
aud[25709]=16'h3243;
aud[25710]=16'h3235;
aud[25711]=16'h3228;
aud[25712]=16'h321b;
aud[25713]=16'h320d;
aud[25714]=16'h3200;
aud[25715]=16'h31f3;
aud[25716]=16'h31e5;
aud[25717]=16'h31d8;
aud[25718]=16'h31ca;
aud[25719]=16'h31bd;
aud[25720]=16'h31af;
aud[25721]=16'h31a2;
aud[25722]=16'h3194;
aud[25723]=16'h3187;
aud[25724]=16'h3179;
aud[25725]=16'h316b;
aud[25726]=16'h315e;
aud[25727]=16'h3150;
aud[25728]=16'h3142;
aud[25729]=16'h3135;
aud[25730]=16'h3127;
aud[25731]=16'h3119;
aud[25732]=16'h310b;
aud[25733]=16'h30fe;
aud[25734]=16'h30f0;
aud[25735]=16'h30e2;
aud[25736]=16'h30d4;
aud[25737]=16'h30c6;
aud[25738]=16'h30b8;
aud[25739]=16'h30aa;
aud[25740]=16'h309d;
aud[25741]=16'h308f;
aud[25742]=16'h3081;
aud[25743]=16'h3073;
aud[25744]=16'h3065;
aud[25745]=16'h3057;
aud[25746]=16'h3048;
aud[25747]=16'h303a;
aud[25748]=16'h302c;
aud[25749]=16'h301e;
aud[25750]=16'h3010;
aud[25751]=16'h3002;
aud[25752]=16'h2ff4;
aud[25753]=16'h2fe5;
aud[25754]=16'h2fd7;
aud[25755]=16'h2fc9;
aud[25756]=16'h2fbb;
aud[25757]=16'h2fac;
aud[25758]=16'h2f9e;
aud[25759]=16'h2f90;
aud[25760]=16'h2f81;
aud[25761]=16'h2f73;
aud[25762]=16'h2f65;
aud[25763]=16'h2f56;
aud[25764]=16'h2f48;
aud[25765]=16'h2f39;
aud[25766]=16'h2f2b;
aud[25767]=16'h2f1c;
aud[25768]=16'h2f0e;
aud[25769]=16'h2eff;
aud[25770]=16'h2ef1;
aud[25771]=16'h2ee2;
aud[25772]=16'h2ed3;
aud[25773]=16'h2ec5;
aud[25774]=16'h2eb6;
aud[25775]=16'h2ea7;
aud[25776]=16'h2e99;
aud[25777]=16'h2e8a;
aud[25778]=16'h2e7b;
aud[25779]=16'h2e6d;
aud[25780]=16'h2e5e;
aud[25781]=16'h2e4f;
aud[25782]=16'h2e40;
aud[25783]=16'h2e31;
aud[25784]=16'h2e22;
aud[25785]=16'h2e14;
aud[25786]=16'h2e05;
aud[25787]=16'h2df6;
aud[25788]=16'h2de7;
aud[25789]=16'h2dd8;
aud[25790]=16'h2dc9;
aud[25791]=16'h2dba;
aud[25792]=16'h2dab;
aud[25793]=16'h2d9c;
aud[25794]=16'h2d8d;
aud[25795]=16'h2d7e;
aud[25796]=16'h2d6f;
aud[25797]=16'h2d60;
aud[25798]=16'h2d50;
aud[25799]=16'h2d41;
aud[25800]=16'h2d32;
aud[25801]=16'h2d23;
aud[25802]=16'h2d14;
aud[25803]=16'h2d04;
aud[25804]=16'h2cf5;
aud[25805]=16'h2ce6;
aud[25806]=16'h2cd7;
aud[25807]=16'h2cc7;
aud[25808]=16'h2cb8;
aud[25809]=16'h2ca9;
aud[25810]=16'h2c99;
aud[25811]=16'h2c8a;
aud[25812]=16'h2c7a;
aud[25813]=16'h2c6b;
aud[25814]=16'h2c5c;
aud[25815]=16'h2c4c;
aud[25816]=16'h2c3d;
aud[25817]=16'h2c2d;
aud[25818]=16'h2c1e;
aud[25819]=16'h2c0e;
aud[25820]=16'h2bfe;
aud[25821]=16'h2bef;
aud[25822]=16'h2bdf;
aud[25823]=16'h2bd0;
aud[25824]=16'h2bc0;
aud[25825]=16'h2bb0;
aud[25826]=16'h2ba1;
aud[25827]=16'h2b91;
aud[25828]=16'h2b81;
aud[25829]=16'h2b71;
aud[25830]=16'h2b62;
aud[25831]=16'h2b52;
aud[25832]=16'h2b42;
aud[25833]=16'h2b32;
aud[25834]=16'h2b22;
aud[25835]=16'h2b13;
aud[25836]=16'h2b03;
aud[25837]=16'h2af3;
aud[25838]=16'h2ae3;
aud[25839]=16'h2ad3;
aud[25840]=16'h2ac3;
aud[25841]=16'h2ab3;
aud[25842]=16'h2aa3;
aud[25843]=16'h2a93;
aud[25844]=16'h2a83;
aud[25845]=16'h2a73;
aud[25846]=16'h2a63;
aud[25847]=16'h2a53;
aud[25848]=16'h2a43;
aud[25849]=16'h2a33;
aud[25850]=16'h2a23;
aud[25851]=16'h2a12;
aud[25852]=16'h2a02;
aud[25853]=16'h29f2;
aud[25854]=16'h29e2;
aud[25855]=16'h29d2;
aud[25856]=16'h29c1;
aud[25857]=16'h29b1;
aud[25858]=16'h29a1;
aud[25859]=16'h2991;
aud[25860]=16'h2980;
aud[25861]=16'h2970;
aud[25862]=16'h2960;
aud[25863]=16'h294f;
aud[25864]=16'h293f;
aud[25865]=16'h292e;
aud[25866]=16'h291e;
aud[25867]=16'h290e;
aud[25868]=16'h28fd;
aud[25869]=16'h28ed;
aud[25870]=16'h28dc;
aud[25871]=16'h28cc;
aud[25872]=16'h28bb;
aud[25873]=16'h28aa;
aud[25874]=16'h289a;
aud[25875]=16'h2889;
aud[25876]=16'h2879;
aud[25877]=16'h2868;
aud[25878]=16'h2857;
aud[25879]=16'h2847;
aud[25880]=16'h2836;
aud[25881]=16'h2825;
aud[25882]=16'h2815;
aud[25883]=16'h2804;
aud[25884]=16'h27f3;
aud[25885]=16'h27e2;
aud[25886]=16'h27d2;
aud[25887]=16'h27c1;
aud[25888]=16'h27b0;
aud[25889]=16'h279f;
aud[25890]=16'h278e;
aud[25891]=16'h277e;
aud[25892]=16'h276d;
aud[25893]=16'h275c;
aud[25894]=16'h274b;
aud[25895]=16'h273a;
aud[25896]=16'h2729;
aud[25897]=16'h2718;
aud[25898]=16'h2707;
aud[25899]=16'h26f6;
aud[25900]=16'h26e5;
aud[25901]=16'h26d4;
aud[25902]=16'h26c3;
aud[25903]=16'h26b2;
aud[25904]=16'h26a1;
aud[25905]=16'h2690;
aud[25906]=16'h267e;
aud[25907]=16'h266d;
aud[25908]=16'h265c;
aud[25909]=16'h264b;
aud[25910]=16'h263a;
aud[25911]=16'h2629;
aud[25912]=16'h2617;
aud[25913]=16'h2606;
aud[25914]=16'h25f5;
aud[25915]=16'h25e4;
aud[25916]=16'h25d2;
aud[25917]=16'h25c1;
aud[25918]=16'h25b0;
aud[25919]=16'h259e;
aud[25920]=16'h258d;
aud[25921]=16'h257c;
aud[25922]=16'h256a;
aud[25923]=16'h2559;
aud[25924]=16'h2547;
aud[25925]=16'h2536;
aud[25926]=16'h2524;
aud[25927]=16'h2513;
aud[25928]=16'h2501;
aud[25929]=16'h24f0;
aud[25930]=16'h24de;
aud[25931]=16'h24cd;
aud[25932]=16'h24bb;
aud[25933]=16'h24aa;
aud[25934]=16'h2498;
aud[25935]=16'h2487;
aud[25936]=16'h2475;
aud[25937]=16'h2463;
aud[25938]=16'h2452;
aud[25939]=16'h2440;
aud[25940]=16'h242e;
aud[25941]=16'h241d;
aud[25942]=16'h240b;
aud[25943]=16'h23f9;
aud[25944]=16'h23e7;
aud[25945]=16'h23d6;
aud[25946]=16'h23c4;
aud[25947]=16'h23b2;
aud[25948]=16'h23a0;
aud[25949]=16'h238e;
aud[25950]=16'h237d;
aud[25951]=16'h236b;
aud[25952]=16'h2359;
aud[25953]=16'h2347;
aud[25954]=16'h2335;
aud[25955]=16'h2323;
aud[25956]=16'h2311;
aud[25957]=16'h22ff;
aud[25958]=16'h22ed;
aud[25959]=16'h22db;
aud[25960]=16'h22c9;
aud[25961]=16'h22b7;
aud[25962]=16'h22a5;
aud[25963]=16'h2293;
aud[25964]=16'h2281;
aud[25965]=16'h226f;
aud[25966]=16'h225d;
aud[25967]=16'h224b;
aud[25968]=16'h2239;
aud[25969]=16'h2227;
aud[25970]=16'h2215;
aud[25971]=16'h2202;
aud[25972]=16'h21f0;
aud[25973]=16'h21de;
aud[25974]=16'h21cc;
aud[25975]=16'h21ba;
aud[25976]=16'h21a7;
aud[25977]=16'h2195;
aud[25978]=16'h2183;
aud[25979]=16'h2171;
aud[25980]=16'h215e;
aud[25981]=16'h214c;
aud[25982]=16'h213a;
aud[25983]=16'h2127;
aud[25984]=16'h2115;
aud[25985]=16'h2103;
aud[25986]=16'h20f0;
aud[25987]=16'h20de;
aud[25988]=16'h20cb;
aud[25989]=16'h20b9;
aud[25990]=16'h20a7;
aud[25991]=16'h2094;
aud[25992]=16'h2082;
aud[25993]=16'h206f;
aud[25994]=16'h205d;
aud[25995]=16'h204a;
aud[25996]=16'h2038;
aud[25997]=16'h2025;
aud[25998]=16'h2013;
aud[25999]=16'h2000;
aud[26000]=16'h1fed;
aud[26001]=16'h1fdb;
aud[26002]=16'h1fc8;
aud[26003]=16'h1fb6;
aud[26004]=16'h1fa3;
aud[26005]=16'h1f90;
aud[26006]=16'h1f7e;
aud[26007]=16'h1f6b;
aud[26008]=16'h1f58;
aud[26009]=16'h1f46;
aud[26010]=16'h1f33;
aud[26011]=16'h1f20;
aud[26012]=16'h1f0d;
aud[26013]=16'h1efb;
aud[26014]=16'h1ee8;
aud[26015]=16'h1ed5;
aud[26016]=16'h1ec2;
aud[26017]=16'h1eaf;
aud[26018]=16'h1e9d;
aud[26019]=16'h1e8a;
aud[26020]=16'h1e77;
aud[26021]=16'h1e64;
aud[26022]=16'h1e51;
aud[26023]=16'h1e3e;
aud[26024]=16'h1e2b;
aud[26025]=16'h1e18;
aud[26026]=16'h1e06;
aud[26027]=16'h1df3;
aud[26028]=16'h1de0;
aud[26029]=16'h1dcd;
aud[26030]=16'h1dba;
aud[26031]=16'h1da7;
aud[26032]=16'h1d94;
aud[26033]=16'h1d81;
aud[26034]=16'h1d6e;
aud[26035]=16'h1d5b;
aud[26036]=16'h1d47;
aud[26037]=16'h1d34;
aud[26038]=16'h1d21;
aud[26039]=16'h1d0e;
aud[26040]=16'h1cfb;
aud[26041]=16'h1ce8;
aud[26042]=16'h1cd5;
aud[26043]=16'h1cc2;
aud[26044]=16'h1cae;
aud[26045]=16'h1c9b;
aud[26046]=16'h1c88;
aud[26047]=16'h1c75;
aud[26048]=16'h1c62;
aud[26049]=16'h1c4e;
aud[26050]=16'h1c3b;
aud[26051]=16'h1c28;
aud[26052]=16'h1c15;
aud[26053]=16'h1c01;
aud[26054]=16'h1bee;
aud[26055]=16'h1bdb;
aud[26056]=16'h1bc8;
aud[26057]=16'h1bb4;
aud[26058]=16'h1ba1;
aud[26059]=16'h1b8d;
aud[26060]=16'h1b7a;
aud[26061]=16'h1b67;
aud[26062]=16'h1b53;
aud[26063]=16'h1b40;
aud[26064]=16'h1b2d;
aud[26065]=16'h1b19;
aud[26066]=16'h1b06;
aud[26067]=16'h1af2;
aud[26068]=16'h1adf;
aud[26069]=16'h1acb;
aud[26070]=16'h1ab8;
aud[26071]=16'h1aa4;
aud[26072]=16'h1a91;
aud[26073]=16'h1a7d;
aud[26074]=16'h1a6a;
aud[26075]=16'h1a56;
aud[26076]=16'h1a43;
aud[26077]=16'h1a2f;
aud[26078]=16'h1a1c;
aud[26079]=16'h1a08;
aud[26080]=16'h19f4;
aud[26081]=16'h19e1;
aud[26082]=16'h19cd;
aud[26083]=16'h19ba;
aud[26084]=16'h19a6;
aud[26085]=16'h1992;
aud[26086]=16'h197f;
aud[26087]=16'h196b;
aud[26088]=16'h1957;
aud[26089]=16'h1943;
aud[26090]=16'h1930;
aud[26091]=16'h191c;
aud[26092]=16'h1908;
aud[26093]=16'h18f5;
aud[26094]=16'h18e1;
aud[26095]=16'h18cd;
aud[26096]=16'h18b9;
aud[26097]=16'h18a5;
aud[26098]=16'h1892;
aud[26099]=16'h187e;
aud[26100]=16'h186a;
aud[26101]=16'h1856;
aud[26102]=16'h1842;
aud[26103]=16'h182f;
aud[26104]=16'h181b;
aud[26105]=16'h1807;
aud[26106]=16'h17f3;
aud[26107]=16'h17df;
aud[26108]=16'h17cb;
aud[26109]=16'h17b7;
aud[26110]=16'h17a3;
aud[26111]=16'h178f;
aud[26112]=16'h177b;
aud[26113]=16'h1767;
aud[26114]=16'h1753;
aud[26115]=16'h1740;
aud[26116]=16'h172c;
aud[26117]=16'h1718;
aud[26118]=16'h1704;
aud[26119]=16'h16f0;
aud[26120]=16'h16db;
aud[26121]=16'h16c7;
aud[26122]=16'h16b3;
aud[26123]=16'h169f;
aud[26124]=16'h168b;
aud[26125]=16'h1677;
aud[26126]=16'h1663;
aud[26127]=16'h164f;
aud[26128]=16'h163b;
aud[26129]=16'h1627;
aud[26130]=16'h1613;
aud[26131]=16'h15ff;
aud[26132]=16'h15ea;
aud[26133]=16'h15d6;
aud[26134]=16'h15c2;
aud[26135]=16'h15ae;
aud[26136]=16'h159a;
aud[26137]=16'h1586;
aud[26138]=16'h1571;
aud[26139]=16'h155d;
aud[26140]=16'h1549;
aud[26141]=16'h1535;
aud[26142]=16'h1520;
aud[26143]=16'h150c;
aud[26144]=16'h14f8;
aud[26145]=16'h14e4;
aud[26146]=16'h14cf;
aud[26147]=16'h14bb;
aud[26148]=16'h14a7;
aud[26149]=16'h1492;
aud[26150]=16'h147e;
aud[26151]=16'h146a;
aud[26152]=16'h1455;
aud[26153]=16'h1441;
aud[26154]=16'h142d;
aud[26155]=16'h1418;
aud[26156]=16'h1404;
aud[26157]=16'h13f0;
aud[26158]=16'h13db;
aud[26159]=16'h13c7;
aud[26160]=16'h13b3;
aud[26161]=16'h139e;
aud[26162]=16'h138a;
aud[26163]=16'h1375;
aud[26164]=16'h1361;
aud[26165]=16'h134c;
aud[26166]=16'h1338;
aud[26167]=16'h1323;
aud[26168]=16'h130f;
aud[26169]=16'h12fb;
aud[26170]=16'h12e6;
aud[26171]=16'h12d2;
aud[26172]=16'h12bd;
aud[26173]=16'h12a9;
aud[26174]=16'h1294;
aud[26175]=16'h127f;
aud[26176]=16'h126b;
aud[26177]=16'h1256;
aud[26178]=16'h1242;
aud[26179]=16'h122d;
aud[26180]=16'h1219;
aud[26181]=16'h1204;
aud[26182]=16'h11f0;
aud[26183]=16'h11db;
aud[26184]=16'h11c6;
aud[26185]=16'h11b2;
aud[26186]=16'h119d;
aud[26187]=16'h1189;
aud[26188]=16'h1174;
aud[26189]=16'h115f;
aud[26190]=16'h114b;
aud[26191]=16'h1136;
aud[26192]=16'h1121;
aud[26193]=16'h110d;
aud[26194]=16'h10f8;
aud[26195]=16'h10e3;
aud[26196]=16'h10cf;
aud[26197]=16'h10ba;
aud[26198]=16'h10a5;
aud[26199]=16'h1090;
aud[26200]=16'h107c;
aud[26201]=16'h1067;
aud[26202]=16'h1052;
aud[26203]=16'h103e;
aud[26204]=16'h1029;
aud[26205]=16'h1014;
aud[26206]=16'hfff;
aud[26207]=16'hfeb;
aud[26208]=16'hfd6;
aud[26209]=16'hfc1;
aud[26210]=16'hfac;
aud[26211]=16'hf97;
aud[26212]=16'hf83;
aud[26213]=16'hf6e;
aud[26214]=16'hf59;
aud[26215]=16'hf44;
aud[26216]=16'hf2f;
aud[26217]=16'hf1a;
aud[26218]=16'hf06;
aud[26219]=16'hef1;
aud[26220]=16'hedc;
aud[26221]=16'hec7;
aud[26222]=16'heb2;
aud[26223]=16'he9d;
aud[26224]=16'he88;
aud[26225]=16'he74;
aud[26226]=16'he5f;
aud[26227]=16'he4a;
aud[26228]=16'he35;
aud[26229]=16'he20;
aud[26230]=16'he0b;
aud[26231]=16'hdf6;
aud[26232]=16'hde1;
aud[26233]=16'hdcc;
aud[26234]=16'hdb7;
aud[26235]=16'hda2;
aud[26236]=16'hd8d;
aud[26237]=16'hd78;
aud[26238]=16'hd63;
aud[26239]=16'hd4e;
aud[26240]=16'hd39;
aud[26241]=16'hd24;
aud[26242]=16'hd0f;
aud[26243]=16'hcfa;
aud[26244]=16'hce5;
aud[26245]=16'hcd0;
aud[26246]=16'hcbb;
aud[26247]=16'hca6;
aud[26248]=16'hc91;
aud[26249]=16'hc7c;
aud[26250]=16'hc67;
aud[26251]=16'hc52;
aud[26252]=16'hc3d;
aud[26253]=16'hc28;
aud[26254]=16'hc13;
aud[26255]=16'hbfe;
aud[26256]=16'hbe9;
aud[26257]=16'hbd4;
aud[26258]=16'hbbf;
aud[26259]=16'hbaa;
aud[26260]=16'hb95;
aud[26261]=16'hb80;
aud[26262]=16'hb6a;
aud[26263]=16'hb55;
aud[26264]=16'hb40;
aud[26265]=16'hb2b;
aud[26266]=16'hb16;
aud[26267]=16'hb01;
aud[26268]=16'haec;
aud[26269]=16'had7;
aud[26270]=16'hac1;
aud[26271]=16'haac;
aud[26272]=16'ha97;
aud[26273]=16'ha82;
aud[26274]=16'ha6d;
aud[26275]=16'ha58;
aud[26276]=16'ha43;
aud[26277]=16'ha2d;
aud[26278]=16'ha18;
aud[26279]=16'ha03;
aud[26280]=16'h9ee;
aud[26281]=16'h9d9;
aud[26282]=16'h9c3;
aud[26283]=16'h9ae;
aud[26284]=16'h999;
aud[26285]=16'h984;
aud[26286]=16'h96f;
aud[26287]=16'h959;
aud[26288]=16'h944;
aud[26289]=16'h92f;
aud[26290]=16'h91a;
aud[26291]=16'h905;
aud[26292]=16'h8ef;
aud[26293]=16'h8da;
aud[26294]=16'h8c5;
aud[26295]=16'h8b0;
aud[26296]=16'h89a;
aud[26297]=16'h885;
aud[26298]=16'h870;
aud[26299]=16'h85b;
aud[26300]=16'h845;
aud[26301]=16'h830;
aud[26302]=16'h81b;
aud[26303]=16'h805;
aud[26304]=16'h7f0;
aud[26305]=16'h7db;
aud[26306]=16'h7c6;
aud[26307]=16'h7b0;
aud[26308]=16'h79b;
aud[26309]=16'h786;
aud[26310]=16'h770;
aud[26311]=16'h75b;
aud[26312]=16'h746;
aud[26313]=16'h731;
aud[26314]=16'h71b;
aud[26315]=16'h706;
aud[26316]=16'h6f1;
aud[26317]=16'h6db;
aud[26318]=16'h6c6;
aud[26319]=16'h6b1;
aud[26320]=16'h69b;
aud[26321]=16'h686;
aud[26322]=16'h671;
aud[26323]=16'h65b;
aud[26324]=16'h646;
aud[26325]=16'h631;
aud[26326]=16'h61b;
aud[26327]=16'h606;
aud[26328]=16'h5f1;
aud[26329]=16'h5db;
aud[26330]=16'h5c6;
aud[26331]=16'h5b0;
aud[26332]=16'h59b;
aud[26333]=16'h586;
aud[26334]=16'h570;
aud[26335]=16'h55b;
aud[26336]=16'h546;
aud[26337]=16'h530;
aud[26338]=16'h51b;
aud[26339]=16'h505;
aud[26340]=16'h4f0;
aud[26341]=16'h4db;
aud[26342]=16'h4c5;
aud[26343]=16'h4b0;
aud[26344]=16'h49b;
aud[26345]=16'h485;
aud[26346]=16'h470;
aud[26347]=16'h45a;
aud[26348]=16'h445;
aud[26349]=16'h430;
aud[26350]=16'h41a;
aud[26351]=16'h405;
aud[26352]=16'h3ef;
aud[26353]=16'h3da;
aud[26354]=16'h3c5;
aud[26355]=16'h3af;
aud[26356]=16'h39a;
aud[26357]=16'h384;
aud[26358]=16'h36f;
aud[26359]=16'h359;
aud[26360]=16'h344;
aud[26361]=16'h32f;
aud[26362]=16'h319;
aud[26363]=16'h304;
aud[26364]=16'h2ee;
aud[26365]=16'h2d9;
aud[26366]=16'h2c4;
aud[26367]=16'h2ae;
aud[26368]=16'h299;
aud[26369]=16'h283;
aud[26370]=16'h26e;
aud[26371]=16'h258;
aud[26372]=16'h243;
aud[26373]=16'h22e;
aud[26374]=16'h218;
aud[26375]=16'h203;
aud[26376]=16'h1ed;
aud[26377]=16'h1d8;
aud[26378]=16'h1c2;
aud[26379]=16'h1ad;
aud[26380]=16'h197;
aud[26381]=16'h182;
aud[26382]=16'h16d;
aud[26383]=16'h157;
aud[26384]=16'h142;
aud[26385]=16'h12c;
aud[26386]=16'h117;
aud[26387]=16'h101;
aud[26388]=16'hec;
aud[26389]=16'hd6;
aud[26390]=16'hc1;
aud[26391]=16'hac;
aud[26392]=16'h96;
aud[26393]=16'h81;
aud[26394]=16'h6b;
aud[26395]=16'h56;
aud[26396]=16'h40;
aud[26397]=16'h2b;
aud[26398]=16'h15;
aud[26399]=16'h0;
aud[26400]=16'hffeb;
aud[26401]=16'hffd5;
aud[26402]=16'hffc0;
aud[26403]=16'hffaa;
aud[26404]=16'hff95;
aud[26405]=16'hff7f;
aud[26406]=16'hff6a;
aud[26407]=16'hff54;
aud[26408]=16'hff3f;
aud[26409]=16'hff2a;
aud[26410]=16'hff14;
aud[26411]=16'hfeff;
aud[26412]=16'hfee9;
aud[26413]=16'hfed4;
aud[26414]=16'hfebe;
aud[26415]=16'hfea9;
aud[26416]=16'hfe93;
aud[26417]=16'hfe7e;
aud[26418]=16'hfe69;
aud[26419]=16'hfe53;
aud[26420]=16'hfe3e;
aud[26421]=16'hfe28;
aud[26422]=16'hfe13;
aud[26423]=16'hfdfd;
aud[26424]=16'hfde8;
aud[26425]=16'hfdd2;
aud[26426]=16'hfdbd;
aud[26427]=16'hfda8;
aud[26428]=16'hfd92;
aud[26429]=16'hfd7d;
aud[26430]=16'hfd67;
aud[26431]=16'hfd52;
aud[26432]=16'hfd3c;
aud[26433]=16'hfd27;
aud[26434]=16'hfd12;
aud[26435]=16'hfcfc;
aud[26436]=16'hfce7;
aud[26437]=16'hfcd1;
aud[26438]=16'hfcbc;
aud[26439]=16'hfca7;
aud[26440]=16'hfc91;
aud[26441]=16'hfc7c;
aud[26442]=16'hfc66;
aud[26443]=16'hfc51;
aud[26444]=16'hfc3b;
aud[26445]=16'hfc26;
aud[26446]=16'hfc11;
aud[26447]=16'hfbfb;
aud[26448]=16'hfbe6;
aud[26449]=16'hfbd0;
aud[26450]=16'hfbbb;
aud[26451]=16'hfba6;
aud[26452]=16'hfb90;
aud[26453]=16'hfb7b;
aud[26454]=16'hfb65;
aud[26455]=16'hfb50;
aud[26456]=16'hfb3b;
aud[26457]=16'hfb25;
aud[26458]=16'hfb10;
aud[26459]=16'hfafb;
aud[26460]=16'hfae5;
aud[26461]=16'hfad0;
aud[26462]=16'hfaba;
aud[26463]=16'hfaa5;
aud[26464]=16'hfa90;
aud[26465]=16'hfa7a;
aud[26466]=16'hfa65;
aud[26467]=16'hfa50;
aud[26468]=16'hfa3a;
aud[26469]=16'hfa25;
aud[26470]=16'hfa0f;
aud[26471]=16'hf9fa;
aud[26472]=16'hf9e5;
aud[26473]=16'hf9cf;
aud[26474]=16'hf9ba;
aud[26475]=16'hf9a5;
aud[26476]=16'hf98f;
aud[26477]=16'hf97a;
aud[26478]=16'hf965;
aud[26479]=16'hf94f;
aud[26480]=16'hf93a;
aud[26481]=16'hf925;
aud[26482]=16'hf90f;
aud[26483]=16'hf8fa;
aud[26484]=16'hf8e5;
aud[26485]=16'hf8cf;
aud[26486]=16'hf8ba;
aud[26487]=16'hf8a5;
aud[26488]=16'hf890;
aud[26489]=16'hf87a;
aud[26490]=16'hf865;
aud[26491]=16'hf850;
aud[26492]=16'hf83a;
aud[26493]=16'hf825;
aud[26494]=16'hf810;
aud[26495]=16'hf7fb;
aud[26496]=16'hf7e5;
aud[26497]=16'hf7d0;
aud[26498]=16'hf7bb;
aud[26499]=16'hf7a5;
aud[26500]=16'hf790;
aud[26501]=16'hf77b;
aud[26502]=16'hf766;
aud[26503]=16'hf750;
aud[26504]=16'hf73b;
aud[26505]=16'hf726;
aud[26506]=16'hf711;
aud[26507]=16'hf6fb;
aud[26508]=16'hf6e6;
aud[26509]=16'hf6d1;
aud[26510]=16'hf6bc;
aud[26511]=16'hf6a7;
aud[26512]=16'hf691;
aud[26513]=16'hf67c;
aud[26514]=16'hf667;
aud[26515]=16'hf652;
aud[26516]=16'hf63d;
aud[26517]=16'hf627;
aud[26518]=16'hf612;
aud[26519]=16'hf5fd;
aud[26520]=16'hf5e8;
aud[26521]=16'hf5d3;
aud[26522]=16'hf5bd;
aud[26523]=16'hf5a8;
aud[26524]=16'hf593;
aud[26525]=16'hf57e;
aud[26526]=16'hf569;
aud[26527]=16'hf554;
aud[26528]=16'hf53f;
aud[26529]=16'hf529;
aud[26530]=16'hf514;
aud[26531]=16'hf4ff;
aud[26532]=16'hf4ea;
aud[26533]=16'hf4d5;
aud[26534]=16'hf4c0;
aud[26535]=16'hf4ab;
aud[26536]=16'hf496;
aud[26537]=16'hf480;
aud[26538]=16'hf46b;
aud[26539]=16'hf456;
aud[26540]=16'hf441;
aud[26541]=16'hf42c;
aud[26542]=16'hf417;
aud[26543]=16'hf402;
aud[26544]=16'hf3ed;
aud[26545]=16'hf3d8;
aud[26546]=16'hf3c3;
aud[26547]=16'hf3ae;
aud[26548]=16'hf399;
aud[26549]=16'hf384;
aud[26550]=16'hf36f;
aud[26551]=16'hf35a;
aud[26552]=16'hf345;
aud[26553]=16'hf330;
aud[26554]=16'hf31b;
aud[26555]=16'hf306;
aud[26556]=16'hf2f1;
aud[26557]=16'hf2dc;
aud[26558]=16'hf2c7;
aud[26559]=16'hf2b2;
aud[26560]=16'hf29d;
aud[26561]=16'hf288;
aud[26562]=16'hf273;
aud[26563]=16'hf25e;
aud[26564]=16'hf249;
aud[26565]=16'hf234;
aud[26566]=16'hf21f;
aud[26567]=16'hf20a;
aud[26568]=16'hf1f5;
aud[26569]=16'hf1e0;
aud[26570]=16'hf1cb;
aud[26571]=16'hf1b6;
aud[26572]=16'hf1a1;
aud[26573]=16'hf18c;
aud[26574]=16'hf178;
aud[26575]=16'hf163;
aud[26576]=16'hf14e;
aud[26577]=16'hf139;
aud[26578]=16'hf124;
aud[26579]=16'hf10f;
aud[26580]=16'hf0fa;
aud[26581]=16'hf0e6;
aud[26582]=16'hf0d1;
aud[26583]=16'hf0bc;
aud[26584]=16'hf0a7;
aud[26585]=16'hf092;
aud[26586]=16'hf07d;
aud[26587]=16'hf069;
aud[26588]=16'hf054;
aud[26589]=16'hf03f;
aud[26590]=16'hf02a;
aud[26591]=16'hf015;
aud[26592]=16'hf001;
aud[26593]=16'hefec;
aud[26594]=16'hefd7;
aud[26595]=16'hefc2;
aud[26596]=16'hefae;
aud[26597]=16'hef99;
aud[26598]=16'hef84;
aud[26599]=16'hef70;
aud[26600]=16'hef5b;
aud[26601]=16'hef46;
aud[26602]=16'hef31;
aud[26603]=16'hef1d;
aud[26604]=16'hef08;
aud[26605]=16'heef3;
aud[26606]=16'heedf;
aud[26607]=16'heeca;
aud[26608]=16'heeb5;
aud[26609]=16'heea1;
aud[26610]=16'hee8c;
aud[26611]=16'hee77;
aud[26612]=16'hee63;
aud[26613]=16'hee4e;
aud[26614]=16'hee3a;
aud[26615]=16'hee25;
aud[26616]=16'hee10;
aud[26617]=16'hedfc;
aud[26618]=16'hede7;
aud[26619]=16'hedd3;
aud[26620]=16'hedbe;
aud[26621]=16'hedaa;
aud[26622]=16'hed95;
aud[26623]=16'hed81;
aud[26624]=16'hed6c;
aud[26625]=16'hed57;
aud[26626]=16'hed43;
aud[26627]=16'hed2e;
aud[26628]=16'hed1a;
aud[26629]=16'hed05;
aud[26630]=16'hecf1;
aud[26631]=16'hecdd;
aud[26632]=16'hecc8;
aud[26633]=16'hecb4;
aud[26634]=16'hec9f;
aud[26635]=16'hec8b;
aud[26636]=16'hec76;
aud[26637]=16'hec62;
aud[26638]=16'hec4d;
aud[26639]=16'hec39;
aud[26640]=16'hec25;
aud[26641]=16'hec10;
aud[26642]=16'hebfc;
aud[26643]=16'hebe8;
aud[26644]=16'hebd3;
aud[26645]=16'hebbf;
aud[26646]=16'hebab;
aud[26647]=16'heb96;
aud[26648]=16'heb82;
aud[26649]=16'heb6e;
aud[26650]=16'heb59;
aud[26651]=16'heb45;
aud[26652]=16'heb31;
aud[26653]=16'heb1c;
aud[26654]=16'heb08;
aud[26655]=16'heaf4;
aud[26656]=16'heae0;
aud[26657]=16'heacb;
aud[26658]=16'heab7;
aud[26659]=16'heaa3;
aud[26660]=16'hea8f;
aud[26661]=16'hea7a;
aud[26662]=16'hea66;
aud[26663]=16'hea52;
aud[26664]=16'hea3e;
aud[26665]=16'hea2a;
aud[26666]=16'hea16;
aud[26667]=16'hea01;
aud[26668]=16'he9ed;
aud[26669]=16'he9d9;
aud[26670]=16'he9c5;
aud[26671]=16'he9b1;
aud[26672]=16'he99d;
aud[26673]=16'he989;
aud[26674]=16'he975;
aud[26675]=16'he961;
aud[26676]=16'he94d;
aud[26677]=16'he939;
aud[26678]=16'he925;
aud[26679]=16'he910;
aud[26680]=16'he8fc;
aud[26681]=16'he8e8;
aud[26682]=16'he8d4;
aud[26683]=16'he8c0;
aud[26684]=16'he8ad;
aud[26685]=16'he899;
aud[26686]=16'he885;
aud[26687]=16'he871;
aud[26688]=16'he85d;
aud[26689]=16'he849;
aud[26690]=16'he835;
aud[26691]=16'he821;
aud[26692]=16'he80d;
aud[26693]=16'he7f9;
aud[26694]=16'he7e5;
aud[26695]=16'he7d1;
aud[26696]=16'he7be;
aud[26697]=16'he7aa;
aud[26698]=16'he796;
aud[26699]=16'he782;
aud[26700]=16'he76e;
aud[26701]=16'he75b;
aud[26702]=16'he747;
aud[26703]=16'he733;
aud[26704]=16'he71f;
aud[26705]=16'he70b;
aud[26706]=16'he6f8;
aud[26707]=16'he6e4;
aud[26708]=16'he6d0;
aud[26709]=16'he6bd;
aud[26710]=16'he6a9;
aud[26711]=16'he695;
aud[26712]=16'he681;
aud[26713]=16'he66e;
aud[26714]=16'he65a;
aud[26715]=16'he646;
aud[26716]=16'he633;
aud[26717]=16'he61f;
aud[26718]=16'he60c;
aud[26719]=16'he5f8;
aud[26720]=16'he5e4;
aud[26721]=16'he5d1;
aud[26722]=16'he5bd;
aud[26723]=16'he5aa;
aud[26724]=16'he596;
aud[26725]=16'he583;
aud[26726]=16'he56f;
aud[26727]=16'he55c;
aud[26728]=16'he548;
aud[26729]=16'he535;
aud[26730]=16'he521;
aud[26731]=16'he50e;
aud[26732]=16'he4fa;
aud[26733]=16'he4e7;
aud[26734]=16'he4d3;
aud[26735]=16'he4c0;
aud[26736]=16'he4ad;
aud[26737]=16'he499;
aud[26738]=16'he486;
aud[26739]=16'he473;
aud[26740]=16'he45f;
aud[26741]=16'he44c;
aud[26742]=16'he438;
aud[26743]=16'he425;
aud[26744]=16'he412;
aud[26745]=16'he3ff;
aud[26746]=16'he3eb;
aud[26747]=16'he3d8;
aud[26748]=16'he3c5;
aud[26749]=16'he3b2;
aud[26750]=16'he39e;
aud[26751]=16'he38b;
aud[26752]=16'he378;
aud[26753]=16'he365;
aud[26754]=16'he352;
aud[26755]=16'he33e;
aud[26756]=16'he32b;
aud[26757]=16'he318;
aud[26758]=16'he305;
aud[26759]=16'he2f2;
aud[26760]=16'he2df;
aud[26761]=16'he2cc;
aud[26762]=16'he2b9;
aud[26763]=16'he2a5;
aud[26764]=16'he292;
aud[26765]=16'he27f;
aud[26766]=16'he26c;
aud[26767]=16'he259;
aud[26768]=16'he246;
aud[26769]=16'he233;
aud[26770]=16'he220;
aud[26771]=16'he20d;
aud[26772]=16'he1fa;
aud[26773]=16'he1e8;
aud[26774]=16'he1d5;
aud[26775]=16'he1c2;
aud[26776]=16'he1af;
aud[26777]=16'he19c;
aud[26778]=16'he189;
aud[26779]=16'he176;
aud[26780]=16'he163;
aud[26781]=16'he151;
aud[26782]=16'he13e;
aud[26783]=16'he12b;
aud[26784]=16'he118;
aud[26785]=16'he105;
aud[26786]=16'he0f3;
aud[26787]=16'he0e0;
aud[26788]=16'he0cd;
aud[26789]=16'he0ba;
aud[26790]=16'he0a8;
aud[26791]=16'he095;
aud[26792]=16'he082;
aud[26793]=16'he070;
aud[26794]=16'he05d;
aud[26795]=16'he04a;
aud[26796]=16'he038;
aud[26797]=16'he025;
aud[26798]=16'he013;
aud[26799]=16'he000;
aud[26800]=16'hdfed;
aud[26801]=16'hdfdb;
aud[26802]=16'hdfc8;
aud[26803]=16'hdfb6;
aud[26804]=16'hdfa3;
aud[26805]=16'hdf91;
aud[26806]=16'hdf7e;
aud[26807]=16'hdf6c;
aud[26808]=16'hdf59;
aud[26809]=16'hdf47;
aud[26810]=16'hdf35;
aud[26811]=16'hdf22;
aud[26812]=16'hdf10;
aud[26813]=16'hdefd;
aud[26814]=16'hdeeb;
aud[26815]=16'hded9;
aud[26816]=16'hdec6;
aud[26817]=16'hdeb4;
aud[26818]=16'hdea2;
aud[26819]=16'hde8f;
aud[26820]=16'hde7d;
aud[26821]=16'hde6b;
aud[26822]=16'hde59;
aud[26823]=16'hde46;
aud[26824]=16'hde34;
aud[26825]=16'hde22;
aud[26826]=16'hde10;
aud[26827]=16'hddfe;
aud[26828]=16'hddeb;
aud[26829]=16'hddd9;
aud[26830]=16'hddc7;
aud[26831]=16'hddb5;
aud[26832]=16'hdda3;
aud[26833]=16'hdd91;
aud[26834]=16'hdd7f;
aud[26835]=16'hdd6d;
aud[26836]=16'hdd5b;
aud[26837]=16'hdd49;
aud[26838]=16'hdd37;
aud[26839]=16'hdd25;
aud[26840]=16'hdd13;
aud[26841]=16'hdd01;
aud[26842]=16'hdcef;
aud[26843]=16'hdcdd;
aud[26844]=16'hdccb;
aud[26845]=16'hdcb9;
aud[26846]=16'hdca7;
aud[26847]=16'hdc95;
aud[26848]=16'hdc83;
aud[26849]=16'hdc72;
aud[26850]=16'hdc60;
aud[26851]=16'hdc4e;
aud[26852]=16'hdc3c;
aud[26853]=16'hdc2a;
aud[26854]=16'hdc19;
aud[26855]=16'hdc07;
aud[26856]=16'hdbf5;
aud[26857]=16'hdbe3;
aud[26858]=16'hdbd2;
aud[26859]=16'hdbc0;
aud[26860]=16'hdbae;
aud[26861]=16'hdb9d;
aud[26862]=16'hdb8b;
aud[26863]=16'hdb79;
aud[26864]=16'hdb68;
aud[26865]=16'hdb56;
aud[26866]=16'hdb45;
aud[26867]=16'hdb33;
aud[26868]=16'hdb22;
aud[26869]=16'hdb10;
aud[26870]=16'hdaff;
aud[26871]=16'hdaed;
aud[26872]=16'hdadc;
aud[26873]=16'hdaca;
aud[26874]=16'hdab9;
aud[26875]=16'hdaa7;
aud[26876]=16'hda96;
aud[26877]=16'hda84;
aud[26878]=16'hda73;
aud[26879]=16'hda62;
aud[26880]=16'hda50;
aud[26881]=16'hda3f;
aud[26882]=16'hda2e;
aud[26883]=16'hda1c;
aud[26884]=16'hda0b;
aud[26885]=16'hd9fa;
aud[26886]=16'hd9e9;
aud[26887]=16'hd9d7;
aud[26888]=16'hd9c6;
aud[26889]=16'hd9b5;
aud[26890]=16'hd9a4;
aud[26891]=16'hd993;
aud[26892]=16'hd982;
aud[26893]=16'hd970;
aud[26894]=16'hd95f;
aud[26895]=16'hd94e;
aud[26896]=16'hd93d;
aud[26897]=16'hd92c;
aud[26898]=16'hd91b;
aud[26899]=16'hd90a;
aud[26900]=16'hd8f9;
aud[26901]=16'hd8e8;
aud[26902]=16'hd8d7;
aud[26903]=16'hd8c6;
aud[26904]=16'hd8b5;
aud[26905]=16'hd8a4;
aud[26906]=16'hd893;
aud[26907]=16'hd882;
aud[26908]=16'hd872;
aud[26909]=16'hd861;
aud[26910]=16'hd850;
aud[26911]=16'hd83f;
aud[26912]=16'hd82e;
aud[26913]=16'hd81e;
aud[26914]=16'hd80d;
aud[26915]=16'hd7fc;
aud[26916]=16'hd7eb;
aud[26917]=16'hd7db;
aud[26918]=16'hd7ca;
aud[26919]=16'hd7b9;
aud[26920]=16'hd7a9;
aud[26921]=16'hd798;
aud[26922]=16'hd787;
aud[26923]=16'hd777;
aud[26924]=16'hd766;
aud[26925]=16'hd756;
aud[26926]=16'hd745;
aud[26927]=16'hd734;
aud[26928]=16'hd724;
aud[26929]=16'hd713;
aud[26930]=16'hd703;
aud[26931]=16'hd6f2;
aud[26932]=16'hd6e2;
aud[26933]=16'hd6d2;
aud[26934]=16'hd6c1;
aud[26935]=16'hd6b1;
aud[26936]=16'hd6a0;
aud[26937]=16'hd690;
aud[26938]=16'hd680;
aud[26939]=16'hd66f;
aud[26940]=16'hd65f;
aud[26941]=16'hd64f;
aud[26942]=16'hd63f;
aud[26943]=16'hd62e;
aud[26944]=16'hd61e;
aud[26945]=16'hd60e;
aud[26946]=16'hd5fe;
aud[26947]=16'hd5ee;
aud[26948]=16'hd5dd;
aud[26949]=16'hd5cd;
aud[26950]=16'hd5bd;
aud[26951]=16'hd5ad;
aud[26952]=16'hd59d;
aud[26953]=16'hd58d;
aud[26954]=16'hd57d;
aud[26955]=16'hd56d;
aud[26956]=16'hd55d;
aud[26957]=16'hd54d;
aud[26958]=16'hd53d;
aud[26959]=16'hd52d;
aud[26960]=16'hd51d;
aud[26961]=16'hd50d;
aud[26962]=16'hd4fd;
aud[26963]=16'hd4ed;
aud[26964]=16'hd4de;
aud[26965]=16'hd4ce;
aud[26966]=16'hd4be;
aud[26967]=16'hd4ae;
aud[26968]=16'hd49e;
aud[26969]=16'hd48f;
aud[26970]=16'hd47f;
aud[26971]=16'hd46f;
aud[26972]=16'hd45f;
aud[26973]=16'hd450;
aud[26974]=16'hd440;
aud[26975]=16'hd430;
aud[26976]=16'hd421;
aud[26977]=16'hd411;
aud[26978]=16'hd402;
aud[26979]=16'hd3f2;
aud[26980]=16'hd3e2;
aud[26981]=16'hd3d3;
aud[26982]=16'hd3c3;
aud[26983]=16'hd3b4;
aud[26984]=16'hd3a4;
aud[26985]=16'hd395;
aud[26986]=16'hd386;
aud[26987]=16'hd376;
aud[26988]=16'hd367;
aud[26989]=16'hd357;
aud[26990]=16'hd348;
aud[26991]=16'hd339;
aud[26992]=16'hd329;
aud[26993]=16'hd31a;
aud[26994]=16'hd30b;
aud[26995]=16'hd2fc;
aud[26996]=16'hd2ec;
aud[26997]=16'hd2dd;
aud[26998]=16'hd2ce;
aud[26999]=16'hd2bf;
aud[27000]=16'hd2b0;
aud[27001]=16'hd2a0;
aud[27002]=16'hd291;
aud[27003]=16'hd282;
aud[27004]=16'hd273;
aud[27005]=16'hd264;
aud[27006]=16'hd255;
aud[27007]=16'hd246;
aud[27008]=16'hd237;
aud[27009]=16'hd228;
aud[27010]=16'hd219;
aud[27011]=16'hd20a;
aud[27012]=16'hd1fb;
aud[27013]=16'hd1ec;
aud[27014]=16'hd1de;
aud[27015]=16'hd1cf;
aud[27016]=16'hd1c0;
aud[27017]=16'hd1b1;
aud[27018]=16'hd1a2;
aud[27019]=16'hd193;
aud[27020]=16'hd185;
aud[27021]=16'hd176;
aud[27022]=16'hd167;
aud[27023]=16'hd159;
aud[27024]=16'hd14a;
aud[27025]=16'hd13b;
aud[27026]=16'hd12d;
aud[27027]=16'hd11e;
aud[27028]=16'hd10f;
aud[27029]=16'hd101;
aud[27030]=16'hd0f2;
aud[27031]=16'hd0e4;
aud[27032]=16'hd0d5;
aud[27033]=16'hd0c7;
aud[27034]=16'hd0b8;
aud[27035]=16'hd0aa;
aud[27036]=16'hd09b;
aud[27037]=16'hd08d;
aud[27038]=16'hd07f;
aud[27039]=16'hd070;
aud[27040]=16'hd062;
aud[27041]=16'hd054;
aud[27042]=16'hd045;
aud[27043]=16'hd037;
aud[27044]=16'hd029;
aud[27045]=16'hd01b;
aud[27046]=16'hd00c;
aud[27047]=16'hcffe;
aud[27048]=16'hcff0;
aud[27049]=16'hcfe2;
aud[27050]=16'hcfd4;
aud[27051]=16'hcfc6;
aud[27052]=16'hcfb8;
aud[27053]=16'hcfa9;
aud[27054]=16'hcf9b;
aud[27055]=16'hcf8d;
aud[27056]=16'hcf7f;
aud[27057]=16'hcf71;
aud[27058]=16'hcf63;
aud[27059]=16'hcf56;
aud[27060]=16'hcf48;
aud[27061]=16'hcf3a;
aud[27062]=16'hcf2c;
aud[27063]=16'hcf1e;
aud[27064]=16'hcf10;
aud[27065]=16'hcf02;
aud[27066]=16'hcef5;
aud[27067]=16'hcee7;
aud[27068]=16'hced9;
aud[27069]=16'hcecb;
aud[27070]=16'hcebe;
aud[27071]=16'hceb0;
aud[27072]=16'hcea2;
aud[27073]=16'hce95;
aud[27074]=16'hce87;
aud[27075]=16'hce79;
aud[27076]=16'hce6c;
aud[27077]=16'hce5e;
aud[27078]=16'hce51;
aud[27079]=16'hce43;
aud[27080]=16'hce36;
aud[27081]=16'hce28;
aud[27082]=16'hce1b;
aud[27083]=16'hce0d;
aud[27084]=16'hce00;
aud[27085]=16'hcdf3;
aud[27086]=16'hcde5;
aud[27087]=16'hcdd8;
aud[27088]=16'hcdcb;
aud[27089]=16'hcdbd;
aud[27090]=16'hcdb0;
aud[27091]=16'hcda3;
aud[27092]=16'hcd96;
aud[27093]=16'hcd88;
aud[27094]=16'hcd7b;
aud[27095]=16'hcd6e;
aud[27096]=16'hcd61;
aud[27097]=16'hcd54;
aud[27098]=16'hcd47;
aud[27099]=16'hcd3a;
aud[27100]=16'hcd2d;
aud[27101]=16'hcd20;
aud[27102]=16'hcd13;
aud[27103]=16'hcd06;
aud[27104]=16'hccf9;
aud[27105]=16'hccec;
aud[27106]=16'hccdf;
aud[27107]=16'hccd2;
aud[27108]=16'hccc5;
aud[27109]=16'hccb8;
aud[27110]=16'hccab;
aud[27111]=16'hcc9f;
aud[27112]=16'hcc92;
aud[27113]=16'hcc85;
aud[27114]=16'hcc78;
aud[27115]=16'hcc6c;
aud[27116]=16'hcc5f;
aud[27117]=16'hcc52;
aud[27118]=16'hcc46;
aud[27119]=16'hcc39;
aud[27120]=16'hcc2c;
aud[27121]=16'hcc20;
aud[27122]=16'hcc13;
aud[27123]=16'hcc07;
aud[27124]=16'hcbfa;
aud[27125]=16'hcbee;
aud[27126]=16'hcbe1;
aud[27127]=16'hcbd5;
aud[27128]=16'hcbc9;
aud[27129]=16'hcbbc;
aud[27130]=16'hcbb0;
aud[27131]=16'hcba3;
aud[27132]=16'hcb97;
aud[27133]=16'hcb8b;
aud[27134]=16'hcb7f;
aud[27135]=16'hcb72;
aud[27136]=16'hcb66;
aud[27137]=16'hcb5a;
aud[27138]=16'hcb4e;
aud[27139]=16'hcb42;
aud[27140]=16'hcb35;
aud[27141]=16'hcb29;
aud[27142]=16'hcb1d;
aud[27143]=16'hcb11;
aud[27144]=16'hcb05;
aud[27145]=16'hcaf9;
aud[27146]=16'hcaed;
aud[27147]=16'hcae1;
aud[27148]=16'hcad5;
aud[27149]=16'hcac9;
aud[27150]=16'hcabd;
aud[27151]=16'hcab1;
aud[27152]=16'hcaa6;
aud[27153]=16'hca9a;
aud[27154]=16'hca8e;
aud[27155]=16'hca82;
aud[27156]=16'hca76;
aud[27157]=16'hca6b;
aud[27158]=16'hca5f;
aud[27159]=16'hca53;
aud[27160]=16'hca48;
aud[27161]=16'hca3c;
aud[27162]=16'hca30;
aud[27163]=16'hca25;
aud[27164]=16'hca19;
aud[27165]=16'hca0e;
aud[27166]=16'hca02;
aud[27167]=16'hc9f7;
aud[27168]=16'hc9eb;
aud[27169]=16'hc9e0;
aud[27170]=16'hc9d4;
aud[27171]=16'hc9c9;
aud[27172]=16'hc9bd;
aud[27173]=16'hc9b2;
aud[27174]=16'hc9a7;
aud[27175]=16'hc99b;
aud[27176]=16'hc990;
aud[27177]=16'hc985;
aud[27178]=16'hc97a;
aud[27179]=16'hc96e;
aud[27180]=16'hc963;
aud[27181]=16'hc958;
aud[27182]=16'hc94d;
aud[27183]=16'hc942;
aud[27184]=16'hc937;
aud[27185]=16'hc92c;
aud[27186]=16'hc920;
aud[27187]=16'hc915;
aud[27188]=16'hc90a;
aud[27189]=16'hc8ff;
aud[27190]=16'hc8f5;
aud[27191]=16'hc8ea;
aud[27192]=16'hc8df;
aud[27193]=16'hc8d4;
aud[27194]=16'hc8c9;
aud[27195]=16'hc8be;
aud[27196]=16'hc8b3;
aud[27197]=16'hc8a9;
aud[27198]=16'hc89e;
aud[27199]=16'hc893;
aud[27200]=16'hc888;
aud[27201]=16'hc87e;
aud[27202]=16'hc873;
aud[27203]=16'hc868;
aud[27204]=16'hc85e;
aud[27205]=16'hc853;
aud[27206]=16'hc849;
aud[27207]=16'hc83e;
aud[27208]=16'hc834;
aud[27209]=16'hc829;
aud[27210]=16'hc81f;
aud[27211]=16'hc814;
aud[27212]=16'hc80a;
aud[27213]=16'hc7ff;
aud[27214]=16'hc7f5;
aud[27215]=16'hc7eb;
aud[27216]=16'hc7e0;
aud[27217]=16'hc7d6;
aud[27218]=16'hc7cc;
aud[27219]=16'hc7c1;
aud[27220]=16'hc7b7;
aud[27221]=16'hc7ad;
aud[27222]=16'hc7a3;
aud[27223]=16'hc799;
aud[27224]=16'hc78f;
aud[27225]=16'hc785;
aud[27226]=16'hc77a;
aud[27227]=16'hc770;
aud[27228]=16'hc766;
aud[27229]=16'hc75c;
aud[27230]=16'hc752;
aud[27231]=16'hc748;
aud[27232]=16'hc73f;
aud[27233]=16'hc735;
aud[27234]=16'hc72b;
aud[27235]=16'hc721;
aud[27236]=16'hc717;
aud[27237]=16'hc70d;
aud[27238]=16'hc703;
aud[27239]=16'hc6fa;
aud[27240]=16'hc6f0;
aud[27241]=16'hc6e6;
aud[27242]=16'hc6dd;
aud[27243]=16'hc6d3;
aud[27244]=16'hc6c9;
aud[27245]=16'hc6c0;
aud[27246]=16'hc6b6;
aud[27247]=16'hc6ad;
aud[27248]=16'hc6a3;
aud[27249]=16'hc69a;
aud[27250]=16'hc690;
aud[27251]=16'hc687;
aud[27252]=16'hc67d;
aud[27253]=16'hc674;
aud[27254]=16'hc66b;
aud[27255]=16'hc661;
aud[27256]=16'hc658;
aud[27257]=16'hc64f;
aud[27258]=16'hc645;
aud[27259]=16'hc63c;
aud[27260]=16'hc633;
aud[27261]=16'hc62a;
aud[27262]=16'hc620;
aud[27263]=16'hc617;
aud[27264]=16'hc60e;
aud[27265]=16'hc605;
aud[27266]=16'hc5fc;
aud[27267]=16'hc5f3;
aud[27268]=16'hc5ea;
aud[27269]=16'hc5e1;
aud[27270]=16'hc5d8;
aud[27271]=16'hc5cf;
aud[27272]=16'hc5c6;
aud[27273]=16'hc5bd;
aud[27274]=16'hc5b4;
aud[27275]=16'hc5ac;
aud[27276]=16'hc5a3;
aud[27277]=16'hc59a;
aud[27278]=16'hc591;
aud[27279]=16'hc588;
aud[27280]=16'hc580;
aud[27281]=16'hc577;
aud[27282]=16'hc56e;
aud[27283]=16'hc566;
aud[27284]=16'hc55d;
aud[27285]=16'hc555;
aud[27286]=16'hc54c;
aud[27287]=16'hc544;
aud[27288]=16'hc53b;
aud[27289]=16'hc533;
aud[27290]=16'hc52a;
aud[27291]=16'hc522;
aud[27292]=16'hc519;
aud[27293]=16'hc511;
aud[27294]=16'hc509;
aud[27295]=16'hc500;
aud[27296]=16'hc4f8;
aud[27297]=16'hc4f0;
aud[27298]=16'hc4e7;
aud[27299]=16'hc4df;
aud[27300]=16'hc4d7;
aud[27301]=16'hc4cf;
aud[27302]=16'hc4c7;
aud[27303]=16'hc4bf;
aud[27304]=16'hc4b6;
aud[27305]=16'hc4ae;
aud[27306]=16'hc4a6;
aud[27307]=16'hc49e;
aud[27308]=16'hc496;
aud[27309]=16'hc48e;
aud[27310]=16'hc486;
aud[27311]=16'hc47f;
aud[27312]=16'hc477;
aud[27313]=16'hc46f;
aud[27314]=16'hc467;
aud[27315]=16'hc45f;
aud[27316]=16'hc457;
aud[27317]=16'hc450;
aud[27318]=16'hc448;
aud[27319]=16'hc440;
aud[27320]=16'hc439;
aud[27321]=16'hc431;
aud[27322]=16'hc429;
aud[27323]=16'hc422;
aud[27324]=16'hc41a;
aud[27325]=16'hc413;
aud[27326]=16'hc40b;
aud[27327]=16'hc404;
aud[27328]=16'hc3fc;
aud[27329]=16'hc3f5;
aud[27330]=16'hc3ed;
aud[27331]=16'hc3e6;
aud[27332]=16'hc3df;
aud[27333]=16'hc3d7;
aud[27334]=16'hc3d0;
aud[27335]=16'hc3c9;
aud[27336]=16'hc3c1;
aud[27337]=16'hc3ba;
aud[27338]=16'hc3b3;
aud[27339]=16'hc3ac;
aud[27340]=16'hc3a5;
aud[27341]=16'hc39d;
aud[27342]=16'hc396;
aud[27343]=16'hc38f;
aud[27344]=16'hc388;
aud[27345]=16'hc381;
aud[27346]=16'hc37a;
aud[27347]=16'hc373;
aud[27348]=16'hc36c;
aud[27349]=16'hc365;
aud[27350]=16'hc35f;
aud[27351]=16'hc358;
aud[27352]=16'hc351;
aud[27353]=16'hc34a;
aud[27354]=16'hc343;
aud[27355]=16'hc33d;
aud[27356]=16'hc336;
aud[27357]=16'hc32f;
aud[27358]=16'hc329;
aud[27359]=16'hc322;
aud[27360]=16'hc31b;
aud[27361]=16'hc315;
aud[27362]=16'hc30e;
aud[27363]=16'hc308;
aud[27364]=16'hc301;
aud[27365]=16'hc2fb;
aud[27366]=16'hc2f4;
aud[27367]=16'hc2ee;
aud[27368]=16'hc2e7;
aud[27369]=16'hc2e1;
aud[27370]=16'hc2db;
aud[27371]=16'hc2d4;
aud[27372]=16'hc2ce;
aud[27373]=16'hc2c8;
aud[27374]=16'hc2c1;
aud[27375]=16'hc2bb;
aud[27376]=16'hc2b5;
aud[27377]=16'hc2af;
aud[27378]=16'hc2a9;
aud[27379]=16'hc2a3;
aud[27380]=16'hc29d;
aud[27381]=16'hc297;
aud[27382]=16'hc291;
aud[27383]=16'hc28b;
aud[27384]=16'hc285;
aud[27385]=16'hc27f;
aud[27386]=16'hc279;
aud[27387]=16'hc273;
aud[27388]=16'hc26d;
aud[27389]=16'hc267;
aud[27390]=16'hc261;
aud[27391]=16'hc25c;
aud[27392]=16'hc256;
aud[27393]=16'hc250;
aud[27394]=16'hc24a;
aud[27395]=16'hc245;
aud[27396]=16'hc23f;
aud[27397]=16'hc239;
aud[27398]=16'hc234;
aud[27399]=16'hc22e;
aud[27400]=16'hc229;
aud[27401]=16'hc223;
aud[27402]=16'hc21e;
aud[27403]=16'hc218;
aud[27404]=16'hc213;
aud[27405]=16'hc20d;
aud[27406]=16'hc208;
aud[27407]=16'hc203;
aud[27408]=16'hc1fd;
aud[27409]=16'hc1f8;
aud[27410]=16'hc1f3;
aud[27411]=16'hc1ee;
aud[27412]=16'hc1e8;
aud[27413]=16'hc1e3;
aud[27414]=16'hc1de;
aud[27415]=16'hc1d9;
aud[27416]=16'hc1d4;
aud[27417]=16'hc1cf;
aud[27418]=16'hc1ca;
aud[27419]=16'hc1c5;
aud[27420]=16'hc1c0;
aud[27421]=16'hc1bb;
aud[27422]=16'hc1b6;
aud[27423]=16'hc1b1;
aud[27424]=16'hc1ac;
aud[27425]=16'hc1a7;
aud[27426]=16'hc1a2;
aud[27427]=16'hc19e;
aud[27428]=16'hc199;
aud[27429]=16'hc194;
aud[27430]=16'hc18f;
aud[27431]=16'hc18b;
aud[27432]=16'hc186;
aud[27433]=16'hc181;
aud[27434]=16'hc17d;
aud[27435]=16'hc178;
aud[27436]=16'hc174;
aud[27437]=16'hc16f;
aud[27438]=16'hc16b;
aud[27439]=16'hc166;
aud[27440]=16'hc162;
aud[27441]=16'hc15d;
aud[27442]=16'hc159;
aud[27443]=16'hc154;
aud[27444]=16'hc150;
aud[27445]=16'hc14c;
aud[27446]=16'hc147;
aud[27447]=16'hc143;
aud[27448]=16'hc13f;
aud[27449]=16'hc13b;
aud[27450]=16'hc137;
aud[27451]=16'hc133;
aud[27452]=16'hc12e;
aud[27453]=16'hc12a;
aud[27454]=16'hc126;
aud[27455]=16'hc122;
aud[27456]=16'hc11e;
aud[27457]=16'hc11a;
aud[27458]=16'hc116;
aud[27459]=16'hc112;
aud[27460]=16'hc10e;
aud[27461]=16'hc10b;
aud[27462]=16'hc107;
aud[27463]=16'hc103;
aud[27464]=16'hc0ff;
aud[27465]=16'hc0fb;
aud[27466]=16'hc0f8;
aud[27467]=16'hc0f4;
aud[27468]=16'hc0f0;
aud[27469]=16'hc0ed;
aud[27470]=16'hc0e9;
aud[27471]=16'hc0e5;
aud[27472]=16'hc0e2;
aud[27473]=16'hc0de;
aud[27474]=16'hc0db;
aud[27475]=16'hc0d7;
aud[27476]=16'hc0d4;
aud[27477]=16'hc0d0;
aud[27478]=16'hc0cd;
aud[27479]=16'hc0ca;
aud[27480]=16'hc0c6;
aud[27481]=16'hc0c3;
aud[27482]=16'hc0c0;
aud[27483]=16'hc0bd;
aud[27484]=16'hc0b9;
aud[27485]=16'hc0b6;
aud[27486]=16'hc0b3;
aud[27487]=16'hc0b0;
aud[27488]=16'hc0ad;
aud[27489]=16'hc0aa;
aud[27490]=16'hc0a6;
aud[27491]=16'hc0a3;
aud[27492]=16'hc0a0;
aud[27493]=16'hc09d;
aud[27494]=16'hc09b;
aud[27495]=16'hc098;
aud[27496]=16'hc095;
aud[27497]=16'hc092;
aud[27498]=16'hc08f;
aud[27499]=16'hc08c;
aud[27500]=16'hc089;
aud[27501]=16'hc087;
aud[27502]=16'hc084;
aud[27503]=16'hc081;
aud[27504]=16'hc07f;
aud[27505]=16'hc07c;
aud[27506]=16'hc079;
aud[27507]=16'hc077;
aud[27508]=16'hc074;
aud[27509]=16'hc072;
aud[27510]=16'hc06f;
aud[27511]=16'hc06d;
aud[27512]=16'hc06a;
aud[27513]=16'hc068;
aud[27514]=16'hc065;
aud[27515]=16'hc063;
aud[27516]=16'hc061;
aud[27517]=16'hc05e;
aud[27518]=16'hc05c;
aud[27519]=16'hc05a;
aud[27520]=16'hc058;
aud[27521]=16'hc055;
aud[27522]=16'hc053;
aud[27523]=16'hc051;
aud[27524]=16'hc04f;
aud[27525]=16'hc04d;
aud[27526]=16'hc04b;
aud[27527]=16'hc049;
aud[27528]=16'hc047;
aud[27529]=16'hc045;
aud[27530]=16'hc043;
aud[27531]=16'hc041;
aud[27532]=16'hc03f;
aud[27533]=16'hc03d;
aud[27534]=16'hc03b;
aud[27535]=16'hc039;
aud[27536]=16'hc038;
aud[27537]=16'hc036;
aud[27538]=16'hc034;
aud[27539]=16'hc033;
aud[27540]=16'hc031;
aud[27541]=16'hc02f;
aud[27542]=16'hc02e;
aud[27543]=16'hc02c;
aud[27544]=16'hc02a;
aud[27545]=16'hc029;
aud[27546]=16'hc027;
aud[27547]=16'hc026;
aud[27548]=16'hc024;
aud[27549]=16'hc023;
aud[27550]=16'hc022;
aud[27551]=16'hc020;
aud[27552]=16'hc01f;
aud[27553]=16'hc01e;
aud[27554]=16'hc01c;
aud[27555]=16'hc01b;
aud[27556]=16'hc01a;
aud[27557]=16'hc019;
aud[27558]=16'hc018;
aud[27559]=16'hc016;
aud[27560]=16'hc015;
aud[27561]=16'hc014;
aud[27562]=16'hc013;
aud[27563]=16'hc012;
aud[27564]=16'hc011;
aud[27565]=16'hc010;
aud[27566]=16'hc00f;
aud[27567]=16'hc00e;
aud[27568]=16'hc00d;
aud[27569]=16'hc00d;
aud[27570]=16'hc00c;
aud[27571]=16'hc00b;
aud[27572]=16'hc00a;
aud[27573]=16'hc009;
aud[27574]=16'hc009;
aud[27575]=16'hc008;
aud[27576]=16'hc007;
aud[27577]=16'hc007;
aud[27578]=16'hc006;
aud[27579]=16'hc006;
aud[27580]=16'hc005;
aud[27581]=16'hc005;
aud[27582]=16'hc004;
aud[27583]=16'hc004;
aud[27584]=16'hc003;
aud[27585]=16'hc003;
aud[27586]=16'hc002;
aud[27587]=16'hc002;
aud[27588]=16'hc002;
aud[27589]=16'hc001;
aud[27590]=16'hc001;
aud[27591]=16'hc001;
aud[27592]=16'hc001;
aud[27593]=16'hc001;
aud[27594]=16'hc000;
aud[27595]=16'hc000;
aud[27596]=16'hc000;
aud[27597]=16'hc000;
aud[27598]=16'hc000;
aud[27599]=16'hc000;
aud[27600]=16'hc000;
aud[27601]=16'hc000;
aud[27602]=16'hc000;
aud[27603]=16'hc000;
aud[27604]=16'hc000;
aud[27605]=16'hc001;
aud[27606]=16'hc001;
aud[27607]=16'hc001;
aud[27608]=16'hc001;
aud[27609]=16'hc001;
aud[27610]=16'hc002;
aud[27611]=16'hc002;
aud[27612]=16'hc002;
aud[27613]=16'hc003;
aud[27614]=16'hc003;
aud[27615]=16'hc004;
aud[27616]=16'hc004;
aud[27617]=16'hc005;
aud[27618]=16'hc005;
aud[27619]=16'hc006;
aud[27620]=16'hc006;
aud[27621]=16'hc007;
aud[27622]=16'hc007;
aud[27623]=16'hc008;
aud[27624]=16'hc009;
aud[27625]=16'hc009;
aud[27626]=16'hc00a;
aud[27627]=16'hc00b;
aud[27628]=16'hc00c;
aud[27629]=16'hc00d;
aud[27630]=16'hc00d;
aud[27631]=16'hc00e;
aud[27632]=16'hc00f;
aud[27633]=16'hc010;
aud[27634]=16'hc011;
aud[27635]=16'hc012;
aud[27636]=16'hc013;
aud[27637]=16'hc014;
aud[27638]=16'hc015;
aud[27639]=16'hc016;
aud[27640]=16'hc018;
aud[27641]=16'hc019;
aud[27642]=16'hc01a;
aud[27643]=16'hc01b;
aud[27644]=16'hc01c;
aud[27645]=16'hc01e;
aud[27646]=16'hc01f;
aud[27647]=16'hc020;
aud[27648]=16'hc022;
aud[27649]=16'hc023;
aud[27650]=16'hc024;
aud[27651]=16'hc026;
aud[27652]=16'hc027;
aud[27653]=16'hc029;
aud[27654]=16'hc02a;
aud[27655]=16'hc02c;
aud[27656]=16'hc02e;
aud[27657]=16'hc02f;
aud[27658]=16'hc031;
aud[27659]=16'hc033;
aud[27660]=16'hc034;
aud[27661]=16'hc036;
aud[27662]=16'hc038;
aud[27663]=16'hc039;
aud[27664]=16'hc03b;
aud[27665]=16'hc03d;
aud[27666]=16'hc03f;
aud[27667]=16'hc041;
aud[27668]=16'hc043;
aud[27669]=16'hc045;
aud[27670]=16'hc047;
aud[27671]=16'hc049;
aud[27672]=16'hc04b;
aud[27673]=16'hc04d;
aud[27674]=16'hc04f;
aud[27675]=16'hc051;
aud[27676]=16'hc053;
aud[27677]=16'hc055;
aud[27678]=16'hc058;
aud[27679]=16'hc05a;
aud[27680]=16'hc05c;
aud[27681]=16'hc05e;
aud[27682]=16'hc061;
aud[27683]=16'hc063;
aud[27684]=16'hc065;
aud[27685]=16'hc068;
aud[27686]=16'hc06a;
aud[27687]=16'hc06d;
aud[27688]=16'hc06f;
aud[27689]=16'hc072;
aud[27690]=16'hc074;
aud[27691]=16'hc077;
aud[27692]=16'hc079;
aud[27693]=16'hc07c;
aud[27694]=16'hc07f;
aud[27695]=16'hc081;
aud[27696]=16'hc084;
aud[27697]=16'hc087;
aud[27698]=16'hc089;
aud[27699]=16'hc08c;
aud[27700]=16'hc08f;
aud[27701]=16'hc092;
aud[27702]=16'hc095;
aud[27703]=16'hc098;
aud[27704]=16'hc09b;
aud[27705]=16'hc09d;
aud[27706]=16'hc0a0;
aud[27707]=16'hc0a3;
aud[27708]=16'hc0a6;
aud[27709]=16'hc0aa;
aud[27710]=16'hc0ad;
aud[27711]=16'hc0b0;
aud[27712]=16'hc0b3;
aud[27713]=16'hc0b6;
aud[27714]=16'hc0b9;
aud[27715]=16'hc0bd;
aud[27716]=16'hc0c0;
aud[27717]=16'hc0c3;
aud[27718]=16'hc0c6;
aud[27719]=16'hc0ca;
aud[27720]=16'hc0cd;
aud[27721]=16'hc0d0;
aud[27722]=16'hc0d4;
aud[27723]=16'hc0d7;
aud[27724]=16'hc0db;
aud[27725]=16'hc0de;
aud[27726]=16'hc0e2;
aud[27727]=16'hc0e5;
aud[27728]=16'hc0e9;
aud[27729]=16'hc0ed;
aud[27730]=16'hc0f0;
aud[27731]=16'hc0f4;
aud[27732]=16'hc0f8;
aud[27733]=16'hc0fb;
aud[27734]=16'hc0ff;
aud[27735]=16'hc103;
aud[27736]=16'hc107;
aud[27737]=16'hc10b;
aud[27738]=16'hc10e;
aud[27739]=16'hc112;
aud[27740]=16'hc116;
aud[27741]=16'hc11a;
aud[27742]=16'hc11e;
aud[27743]=16'hc122;
aud[27744]=16'hc126;
aud[27745]=16'hc12a;
aud[27746]=16'hc12e;
aud[27747]=16'hc133;
aud[27748]=16'hc137;
aud[27749]=16'hc13b;
aud[27750]=16'hc13f;
aud[27751]=16'hc143;
aud[27752]=16'hc147;
aud[27753]=16'hc14c;
aud[27754]=16'hc150;
aud[27755]=16'hc154;
aud[27756]=16'hc159;
aud[27757]=16'hc15d;
aud[27758]=16'hc162;
aud[27759]=16'hc166;
aud[27760]=16'hc16b;
aud[27761]=16'hc16f;
aud[27762]=16'hc174;
aud[27763]=16'hc178;
aud[27764]=16'hc17d;
aud[27765]=16'hc181;
aud[27766]=16'hc186;
aud[27767]=16'hc18b;
aud[27768]=16'hc18f;
aud[27769]=16'hc194;
aud[27770]=16'hc199;
aud[27771]=16'hc19e;
aud[27772]=16'hc1a2;
aud[27773]=16'hc1a7;
aud[27774]=16'hc1ac;
aud[27775]=16'hc1b1;
aud[27776]=16'hc1b6;
aud[27777]=16'hc1bb;
aud[27778]=16'hc1c0;
aud[27779]=16'hc1c5;
aud[27780]=16'hc1ca;
aud[27781]=16'hc1cf;
aud[27782]=16'hc1d4;
aud[27783]=16'hc1d9;
aud[27784]=16'hc1de;
aud[27785]=16'hc1e3;
aud[27786]=16'hc1e8;
aud[27787]=16'hc1ee;
aud[27788]=16'hc1f3;
aud[27789]=16'hc1f8;
aud[27790]=16'hc1fd;
aud[27791]=16'hc203;
aud[27792]=16'hc208;
aud[27793]=16'hc20d;
aud[27794]=16'hc213;
aud[27795]=16'hc218;
aud[27796]=16'hc21e;
aud[27797]=16'hc223;
aud[27798]=16'hc229;
aud[27799]=16'hc22e;
aud[27800]=16'hc234;
aud[27801]=16'hc239;
aud[27802]=16'hc23f;
aud[27803]=16'hc245;
aud[27804]=16'hc24a;
aud[27805]=16'hc250;
aud[27806]=16'hc256;
aud[27807]=16'hc25c;
aud[27808]=16'hc261;
aud[27809]=16'hc267;
aud[27810]=16'hc26d;
aud[27811]=16'hc273;
aud[27812]=16'hc279;
aud[27813]=16'hc27f;
aud[27814]=16'hc285;
aud[27815]=16'hc28b;
aud[27816]=16'hc291;
aud[27817]=16'hc297;
aud[27818]=16'hc29d;
aud[27819]=16'hc2a3;
aud[27820]=16'hc2a9;
aud[27821]=16'hc2af;
aud[27822]=16'hc2b5;
aud[27823]=16'hc2bb;
aud[27824]=16'hc2c1;
aud[27825]=16'hc2c8;
aud[27826]=16'hc2ce;
aud[27827]=16'hc2d4;
aud[27828]=16'hc2db;
aud[27829]=16'hc2e1;
aud[27830]=16'hc2e7;
aud[27831]=16'hc2ee;
aud[27832]=16'hc2f4;
aud[27833]=16'hc2fb;
aud[27834]=16'hc301;
aud[27835]=16'hc308;
aud[27836]=16'hc30e;
aud[27837]=16'hc315;
aud[27838]=16'hc31b;
aud[27839]=16'hc322;
aud[27840]=16'hc329;
aud[27841]=16'hc32f;
aud[27842]=16'hc336;
aud[27843]=16'hc33d;
aud[27844]=16'hc343;
aud[27845]=16'hc34a;
aud[27846]=16'hc351;
aud[27847]=16'hc358;
aud[27848]=16'hc35f;
aud[27849]=16'hc365;
aud[27850]=16'hc36c;
aud[27851]=16'hc373;
aud[27852]=16'hc37a;
aud[27853]=16'hc381;
aud[27854]=16'hc388;
aud[27855]=16'hc38f;
aud[27856]=16'hc396;
aud[27857]=16'hc39d;
aud[27858]=16'hc3a5;
aud[27859]=16'hc3ac;
aud[27860]=16'hc3b3;
aud[27861]=16'hc3ba;
aud[27862]=16'hc3c1;
aud[27863]=16'hc3c9;
aud[27864]=16'hc3d0;
aud[27865]=16'hc3d7;
aud[27866]=16'hc3df;
aud[27867]=16'hc3e6;
aud[27868]=16'hc3ed;
aud[27869]=16'hc3f5;
aud[27870]=16'hc3fc;
aud[27871]=16'hc404;
aud[27872]=16'hc40b;
aud[27873]=16'hc413;
aud[27874]=16'hc41a;
aud[27875]=16'hc422;
aud[27876]=16'hc429;
aud[27877]=16'hc431;
aud[27878]=16'hc439;
aud[27879]=16'hc440;
aud[27880]=16'hc448;
aud[27881]=16'hc450;
aud[27882]=16'hc457;
aud[27883]=16'hc45f;
aud[27884]=16'hc467;
aud[27885]=16'hc46f;
aud[27886]=16'hc477;
aud[27887]=16'hc47f;
aud[27888]=16'hc486;
aud[27889]=16'hc48e;
aud[27890]=16'hc496;
aud[27891]=16'hc49e;
aud[27892]=16'hc4a6;
aud[27893]=16'hc4ae;
aud[27894]=16'hc4b6;
aud[27895]=16'hc4bf;
aud[27896]=16'hc4c7;
aud[27897]=16'hc4cf;
aud[27898]=16'hc4d7;
aud[27899]=16'hc4df;
aud[27900]=16'hc4e7;
aud[27901]=16'hc4f0;
aud[27902]=16'hc4f8;
aud[27903]=16'hc500;
aud[27904]=16'hc509;
aud[27905]=16'hc511;
aud[27906]=16'hc519;
aud[27907]=16'hc522;
aud[27908]=16'hc52a;
aud[27909]=16'hc533;
aud[27910]=16'hc53b;
aud[27911]=16'hc544;
aud[27912]=16'hc54c;
aud[27913]=16'hc555;
aud[27914]=16'hc55d;
aud[27915]=16'hc566;
aud[27916]=16'hc56e;
aud[27917]=16'hc577;
aud[27918]=16'hc580;
aud[27919]=16'hc588;
aud[27920]=16'hc591;
aud[27921]=16'hc59a;
aud[27922]=16'hc5a3;
aud[27923]=16'hc5ac;
aud[27924]=16'hc5b4;
aud[27925]=16'hc5bd;
aud[27926]=16'hc5c6;
aud[27927]=16'hc5cf;
aud[27928]=16'hc5d8;
aud[27929]=16'hc5e1;
aud[27930]=16'hc5ea;
aud[27931]=16'hc5f3;
aud[27932]=16'hc5fc;
aud[27933]=16'hc605;
aud[27934]=16'hc60e;
aud[27935]=16'hc617;
aud[27936]=16'hc620;
aud[27937]=16'hc62a;
aud[27938]=16'hc633;
aud[27939]=16'hc63c;
aud[27940]=16'hc645;
aud[27941]=16'hc64f;
aud[27942]=16'hc658;
aud[27943]=16'hc661;
aud[27944]=16'hc66b;
aud[27945]=16'hc674;
aud[27946]=16'hc67d;
aud[27947]=16'hc687;
aud[27948]=16'hc690;
aud[27949]=16'hc69a;
aud[27950]=16'hc6a3;
aud[27951]=16'hc6ad;
aud[27952]=16'hc6b6;
aud[27953]=16'hc6c0;
aud[27954]=16'hc6c9;
aud[27955]=16'hc6d3;
aud[27956]=16'hc6dd;
aud[27957]=16'hc6e6;
aud[27958]=16'hc6f0;
aud[27959]=16'hc6fa;
aud[27960]=16'hc703;
aud[27961]=16'hc70d;
aud[27962]=16'hc717;
aud[27963]=16'hc721;
aud[27964]=16'hc72b;
aud[27965]=16'hc735;
aud[27966]=16'hc73f;
aud[27967]=16'hc748;
aud[27968]=16'hc752;
aud[27969]=16'hc75c;
aud[27970]=16'hc766;
aud[27971]=16'hc770;
aud[27972]=16'hc77a;
aud[27973]=16'hc785;
aud[27974]=16'hc78f;
aud[27975]=16'hc799;
aud[27976]=16'hc7a3;
aud[27977]=16'hc7ad;
aud[27978]=16'hc7b7;
aud[27979]=16'hc7c1;
aud[27980]=16'hc7cc;
aud[27981]=16'hc7d6;
aud[27982]=16'hc7e0;
aud[27983]=16'hc7eb;
aud[27984]=16'hc7f5;
aud[27985]=16'hc7ff;
aud[27986]=16'hc80a;
aud[27987]=16'hc814;
aud[27988]=16'hc81f;
aud[27989]=16'hc829;
aud[27990]=16'hc834;
aud[27991]=16'hc83e;
aud[27992]=16'hc849;
aud[27993]=16'hc853;
aud[27994]=16'hc85e;
aud[27995]=16'hc868;
aud[27996]=16'hc873;
aud[27997]=16'hc87e;
aud[27998]=16'hc888;
aud[27999]=16'hc893;
aud[28000]=16'hc89e;
aud[28001]=16'hc8a9;
aud[28002]=16'hc8b3;
aud[28003]=16'hc8be;
aud[28004]=16'hc8c9;
aud[28005]=16'hc8d4;
aud[28006]=16'hc8df;
aud[28007]=16'hc8ea;
aud[28008]=16'hc8f5;
aud[28009]=16'hc8ff;
aud[28010]=16'hc90a;
aud[28011]=16'hc915;
aud[28012]=16'hc920;
aud[28013]=16'hc92c;
aud[28014]=16'hc937;
aud[28015]=16'hc942;
aud[28016]=16'hc94d;
aud[28017]=16'hc958;
aud[28018]=16'hc963;
aud[28019]=16'hc96e;
aud[28020]=16'hc97a;
aud[28021]=16'hc985;
aud[28022]=16'hc990;
aud[28023]=16'hc99b;
aud[28024]=16'hc9a7;
aud[28025]=16'hc9b2;
aud[28026]=16'hc9bd;
aud[28027]=16'hc9c9;
aud[28028]=16'hc9d4;
aud[28029]=16'hc9e0;
aud[28030]=16'hc9eb;
aud[28031]=16'hc9f7;
aud[28032]=16'hca02;
aud[28033]=16'hca0e;
aud[28034]=16'hca19;
aud[28035]=16'hca25;
aud[28036]=16'hca30;
aud[28037]=16'hca3c;
aud[28038]=16'hca48;
aud[28039]=16'hca53;
aud[28040]=16'hca5f;
aud[28041]=16'hca6b;
aud[28042]=16'hca76;
aud[28043]=16'hca82;
aud[28044]=16'hca8e;
aud[28045]=16'hca9a;
aud[28046]=16'hcaa6;
aud[28047]=16'hcab1;
aud[28048]=16'hcabd;
aud[28049]=16'hcac9;
aud[28050]=16'hcad5;
aud[28051]=16'hcae1;
aud[28052]=16'hcaed;
aud[28053]=16'hcaf9;
aud[28054]=16'hcb05;
aud[28055]=16'hcb11;
aud[28056]=16'hcb1d;
aud[28057]=16'hcb29;
aud[28058]=16'hcb35;
aud[28059]=16'hcb42;
aud[28060]=16'hcb4e;
aud[28061]=16'hcb5a;
aud[28062]=16'hcb66;
aud[28063]=16'hcb72;
aud[28064]=16'hcb7f;
aud[28065]=16'hcb8b;
aud[28066]=16'hcb97;
aud[28067]=16'hcba3;
aud[28068]=16'hcbb0;
aud[28069]=16'hcbbc;
aud[28070]=16'hcbc9;
aud[28071]=16'hcbd5;
aud[28072]=16'hcbe1;
aud[28073]=16'hcbee;
aud[28074]=16'hcbfa;
aud[28075]=16'hcc07;
aud[28076]=16'hcc13;
aud[28077]=16'hcc20;
aud[28078]=16'hcc2c;
aud[28079]=16'hcc39;
aud[28080]=16'hcc46;
aud[28081]=16'hcc52;
aud[28082]=16'hcc5f;
aud[28083]=16'hcc6c;
aud[28084]=16'hcc78;
aud[28085]=16'hcc85;
aud[28086]=16'hcc92;
aud[28087]=16'hcc9f;
aud[28088]=16'hccab;
aud[28089]=16'hccb8;
aud[28090]=16'hccc5;
aud[28091]=16'hccd2;
aud[28092]=16'hccdf;
aud[28093]=16'hccec;
aud[28094]=16'hccf9;
aud[28095]=16'hcd06;
aud[28096]=16'hcd13;
aud[28097]=16'hcd20;
aud[28098]=16'hcd2d;
aud[28099]=16'hcd3a;
aud[28100]=16'hcd47;
aud[28101]=16'hcd54;
aud[28102]=16'hcd61;
aud[28103]=16'hcd6e;
aud[28104]=16'hcd7b;
aud[28105]=16'hcd88;
aud[28106]=16'hcd96;
aud[28107]=16'hcda3;
aud[28108]=16'hcdb0;
aud[28109]=16'hcdbd;
aud[28110]=16'hcdcb;
aud[28111]=16'hcdd8;
aud[28112]=16'hcde5;
aud[28113]=16'hcdf3;
aud[28114]=16'hce00;
aud[28115]=16'hce0d;
aud[28116]=16'hce1b;
aud[28117]=16'hce28;
aud[28118]=16'hce36;
aud[28119]=16'hce43;
aud[28120]=16'hce51;
aud[28121]=16'hce5e;
aud[28122]=16'hce6c;
aud[28123]=16'hce79;
aud[28124]=16'hce87;
aud[28125]=16'hce95;
aud[28126]=16'hcea2;
aud[28127]=16'hceb0;
aud[28128]=16'hcebe;
aud[28129]=16'hcecb;
aud[28130]=16'hced9;
aud[28131]=16'hcee7;
aud[28132]=16'hcef5;
aud[28133]=16'hcf02;
aud[28134]=16'hcf10;
aud[28135]=16'hcf1e;
aud[28136]=16'hcf2c;
aud[28137]=16'hcf3a;
aud[28138]=16'hcf48;
aud[28139]=16'hcf56;
aud[28140]=16'hcf63;
aud[28141]=16'hcf71;
aud[28142]=16'hcf7f;
aud[28143]=16'hcf8d;
aud[28144]=16'hcf9b;
aud[28145]=16'hcfa9;
aud[28146]=16'hcfb8;
aud[28147]=16'hcfc6;
aud[28148]=16'hcfd4;
aud[28149]=16'hcfe2;
aud[28150]=16'hcff0;
aud[28151]=16'hcffe;
aud[28152]=16'hd00c;
aud[28153]=16'hd01b;
aud[28154]=16'hd029;
aud[28155]=16'hd037;
aud[28156]=16'hd045;
aud[28157]=16'hd054;
aud[28158]=16'hd062;
aud[28159]=16'hd070;
aud[28160]=16'hd07f;
aud[28161]=16'hd08d;
aud[28162]=16'hd09b;
aud[28163]=16'hd0aa;
aud[28164]=16'hd0b8;
aud[28165]=16'hd0c7;
aud[28166]=16'hd0d5;
aud[28167]=16'hd0e4;
aud[28168]=16'hd0f2;
aud[28169]=16'hd101;
aud[28170]=16'hd10f;
aud[28171]=16'hd11e;
aud[28172]=16'hd12d;
aud[28173]=16'hd13b;
aud[28174]=16'hd14a;
aud[28175]=16'hd159;
aud[28176]=16'hd167;
aud[28177]=16'hd176;
aud[28178]=16'hd185;
aud[28179]=16'hd193;
aud[28180]=16'hd1a2;
aud[28181]=16'hd1b1;
aud[28182]=16'hd1c0;
aud[28183]=16'hd1cf;
aud[28184]=16'hd1de;
aud[28185]=16'hd1ec;
aud[28186]=16'hd1fb;
aud[28187]=16'hd20a;
aud[28188]=16'hd219;
aud[28189]=16'hd228;
aud[28190]=16'hd237;
aud[28191]=16'hd246;
aud[28192]=16'hd255;
aud[28193]=16'hd264;
aud[28194]=16'hd273;
aud[28195]=16'hd282;
aud[28196]=16'hd291;
aud[28197]=16'hd2a0;
aud[28198]=16'hd2b0;
aud[28199]=16'hd2bf;
aud[28200]=16'hd2ce;
aud[28201]=16'hd2dd;
aud[28202]=16'hd2ec;
aud[28203]=16'hd2fc;
aud[28204]=16'hd30b;
aud[28205]=16'hd31a;
aud[28206]=16'hd329;
aud[28207]=16'hd339;
aud[28208]=16'hd348;
aud[28209]=16'hd357;
aud[28210]=16'hd367;
aud[28211]=16'hd376;
aud[28212]=16'hd386;
aud[28213]=16'hd395;
aud[28214]=16'hd3a4;
aud[28215]=16'hd3b4;
aud[28216]=16'hd3c3;
aud[28217]=16'hd3d3;
aud[28218]=16'hd3e2;
aud[28219]=16'hd3f2;
aud[28220]=16'hd402;
aud[28221]=16'hd411;
aud[28222]=16'hd421;
aud[28223]=16'hd430;
aud[28224]=16'hd440;
aud[28225]=16'hd450;
aud[28226]=16'hd45f;
aud[28227]=16'hd46f;
aud[28228]=16'hd47f;
aud[28229]=16'hd48f;
aud[28230]=16'hd49e;
aud[28231]=16'hd4ae;
aud[28232]=16'hd4be;
aud[28233]=16'hd4ce;
aud[28234]=16'hd4de;
aud[28235]=16'hd4ed;
aud[28236]=16'hd4fd;
aud[28237]=16'hd50d;
aud[28238]=16'hd51d;
aud[28239]=16'hd52d;
aud[28240]=16'hd53d;
aud[28241]=16'hd54d;
aud[28242]=16'hd55d;
aud[28243]=16'hd56d;
aud[28244]=16'hd57d;
aud[28245]=16'hd58d;
aud[28246]=16'hd59d;
aud[28247]=16'hd5ad;
aud[28248]=16'hd5bd;
aud[28249]=16'hd5cd;
aud[28250]=16'hd5dd;
aud[28251]=16'hd5ee;
aud[28252]=16'hd5fe;
aud[28253]=16'hd60e;
aud[28254]=16'hd61e;
aud[28255]=16'hd62e;
aud[28256]=16'hd63f;
aud[28257]=16'hd64f;
aud[28258]=16'hd65f;
aud[28259]=16'hd66f;
aud[28260]=16'hd680;
aud[28261]=16'hd690;
aud[28262]=16'hd6a0;
aud[28263]=16'hd6b1;
aud[28264]=16'hd6c1;
aud[28265]=16'hd6d2;
aud[28266]=16'hd6e2;
aud[28267]=16'hd6f2;
aud[28268]=16'hd703;
aud[28269]=16'hd713;
aud[28270]=16'hd724;
aud[28271]=16'hd734;
aud[28272]=16'hd745;
aud[28273]=16'hd756;
aud[28274]=16'hd766;
aud[28275]=16'hd777;
aud[28276]=16'hd787;
aud[28277]=16'hd798;
aud[28278]=16'hd7a9;
aud[28279]=16'hd7b9;
aud[28280]=16'hd7ca;
aud[28281]=16'hd7db;
aud[28282]=16'hd7eb;
aud[28283]=16'hd7fc;
aud[28284]=16'hd80d;
aud[28285]=16'hd81e;
aud[28286]=16'hd82e;
aud[28287]=16'hd83f;
aud[28288]=16'hd850;
aud[28289]=16'hd861;
aud[28290]=16'hd872;
aud[28291]=16'hd882;
aud[28292]=16'hd893;
aud[28293]=16'hd8a4;
aud[28294]=16'hd8b5;
aud[28295]=16'hd8c6;
aud[28296]=16'hd8d7;
aud[28297]=16'hd8e8;
aud[28298]=16'hd8f9;
aud[28299]=16'hd90a;
aud[28300]=16'hd91b;
aud[28301]=16'hd92c;
aud[28302]=16'hd93d;
aud[28303]=16'hd94e;
aud[28304]=16'hd95f;
aud[28305]=16'hd970;
aud[28306]=16'hd982;
aud[28307]=16'hd993;
aud[28308]=16'hd9a4;
aud[28309]=16'hd9b5;
aud[28310]=16'hd9c6;
aud[28311]=16'hd9d7;
aud[28312]=16'hd9e9;
aud[28313]=16'hd9fa;
aud[28314]=16'hda0b;
aud[28315]=16'hda1c;
aud[28316]=16'hda2e;
aud[28317]=16'hda3f;
aud[28318]=16'hda50;
aud[28319]=16'hda62;
aud[28320]=16'hda73;
aud[28321]=16'hda84;
aud[28322]=16'hda96;
aud[28323]=16'hdaa7;
aud[28324]=16'hdab9;
aud[28325]=16'hdaca;
aud[28326]=16'hdadc;
aud[28327]=16'hdaed;
aud[28328]=16'hdaff;
aud[28329]=16'hdb10;
aud[28330]=16'hdb22;
aud[28331]=16'hdb33;
aud[28332]=16'hdb45;
aud[28333]=16'hdb56;
aud[28334]=16'hdb68;
aud[28335]=16'hdb79;
aud[28336]=16'hdb8b;
aud[28337]=16'hdb9d;
aud[28338]=16'hdbae;
aud[28339]=16'hdbc0;
aud[28340]=16'hdbd2;
aud[28341]=16'hdbe3;
aud[28342]=16'hdbf5;
aud[28343]=16'hdc07;
aud[28344]=16'hdc19;
aud[28345]=16'hdc2a;
aud[28346]=16'hdc3c;
aud[28347]=16'hdc4e;
aud[28348]=16'hdc60;
aud[28349]=16'hdc72;
aud[28350]=16'hdc83;
aud[28351]=16'hdc95;
aud[28352]=16'hdca7;
aud[28353]=16'hdcb9;
aud[28354]=16'hdccb;
aud[28355]=16'hdcdd;
aud[28356]=16'hdcef;
aud[28357]=16'hdd01;
aud[28358]=16'hdd13;
aud[28359]=16'hdd25;
aud[28360]=16'hdd37;
aud[28361]=16'hdd49;
aud[28362]=16'hdd5b;
aud[28363]=16'hdd6d;
aud[28364]=16'hdd7f;
aud[28365]=16'hdd91;
aud[28366]=16'hdda3;
aud[28367]=16'hddb5;
aud[28368]=16'hddc7;
aud[28369]=16'hddd9;
aud[28370]=16'hddeb;
aud[28371]=16'hddfe;
aud[28372]=16'hde10;
aud[28373]=16'hde22;
aud[28374]=16'hde34;
aud[28375]=16'hde46;
aud[28376]=16'hde59;
aud[28377]=16'hde6b;
aud[28378]=16'hde7d;
aud[28379]=16'hde8f;
aud[28380]=16'hdea2;
aud[28381]=16'hdeb4;
aud[28382]=16'hdec6;
aud[28383]=16'hded9;
aud[28384]=16'hdeeb;
aud[28385]=16'hdefd;
aud[28386]=16'hdf10;
aud[28387]=16'hdf22;
aud[28388]=16'hdf35;
aud[28389]=16'hdf47;
aud[28390]=16'hdf59;
aud[28391]=16'hdf6c;
aud[28392]=16'hdf7e;
aud[28393]=16'hdf91;
aud[28394]=16'hdfa3;
aud[28395]=16'hdfb6;
aud[28396]=16'hdfc8;
aud[28397]=16'hdfdb;
aud[28398]=16'hdfed;
aud[28399]=16'he000;
aud[28400]=16'he013;
aud[28401]=16'he025;
aud[28402]=16'he038;
aud[28403]=16'he04a;
aud[28404]=16'he05d;
aud[28405]=16'he070;
aud[28406]=16'he082;
aud[28407]=16'he095;
aud[28408]=16'he0a8;
aud[28409]=16'he0ba;
aud[28410]=16'he0cd;
aud[28411]=16'he0e0;
aud[28412]=16'he0f3;
aud[28413]=16'he105;
aud[28414]=16'he118;
aud[28415]=16'he12b;
aud[28416]=16'he13e;
aud[28417]=16'he151;
aud[28418]=16'he163;
aud[28419]=16'he176;
aud[28420]=16'he189;
aud[28421]=16'he19c;
aud[28422]=16'he1af;
aud[28423]=16'he1c2;
aud[28424]=16'he1d5;
aud[28425]=16'he1e8;
aud[28426]=16'he1fa;
aud[28427]=16'he20d;
aud[28428]=16'he220;
aud[28429]=16'he233;
aud[28430]=16'he246;
aud[28431]=16'he259;
aud[28432]=16'he26c;
aud[28433]=16'he27f;
aud[28434]=16'he292;
aud[28435]=16'he2a5;
aud[28436]=16'he2b9;
aud[28437]=16'he2cc;
aud[28438]=16'he2df;
aud[28439]=16'he2f2;
aud[28440]=16'he305;
aud[28441]=16'he318;
aud[28442]=16'he32b;
aud[28443]=16'he33e;
aud[28444]=16'he352;
aud[28445]=16'he365;
aud[28446]=16'he378;
aud[28447]=16'he38b;
aud[28448]=16'he39e;
aud[28449]=16'he3b2;
aud[28450]=16'he3c5;
aud[28451]=16'he3d8;
aud[28452]=16'he3eb;
aud[28453]=16'he3ff;
aud[28454]=16'he412;
aud[28455]=16'he425;
aud[28456]=16'he438;
aud[28457]=16'he44c;
aud[28458]=16'he45f;
aud[28459]=16'he473;
aud[28460]=16'he486;
aud[28461]=16'he499;
aud[28462]=16'he4ad;
aud[28463]=16'he4c0;
aud[28464]=16'he4d3;
aud[28465]=16'he4e7;
aud[28466]=16'he4fa;
aud[28467]=16'he50e;
aud[28468]=16'he521;
aud[28469]=16'he535;
aud[28470]=16'he548;
aud[28471]=16'he55c;
aud[28472]=16'he56f;
aud[28473]=16'he583;
aud[28474]=16'he596;
aud[28475]=16'he5aa;
aud[28476]=16'he5bd;
aud[28477]=16'he5d1;
aud[28478]=16'he5e4;
aud[28479]=16'he5f8;
aud[28480]=16'he60c;
aud[28481]=16'he61f;
aud[28482]=16'he633;
aud[28483]=16'he646;
aud[28484]=16'he65a;
aud[28485]=16'he66e;
aud[28486]=16'he681;
aud[28487]=16'he695;
aud[28488]=16'he6a9;
aud[28489]=16'he6bd;
aud[28490]=16'he6d0;
aud[28491]=16'he6e4;
aud[28492]=16'he6f8;
aud[28493]=16'he70b;
aud[28494]=16'he71f;
aud[28495]=16'he733;
aud[28496]=16'he747;
aud[28497]=16'he75b;
aud[28498]=16'he76e;
aud[28499]=16'he782;
aud[28500]=16'he796;
aud[28501]=16'he7aa;
aud[28502]=16'he7be;
aud[28503]=16'he7d1;
aud[28504]=16'he7e5;
aud[28505]=16'he7f9;
aud[28506]=16'he80d;
aud[28507]=16'he821;
aud[28508]=16'he835;
aud[28509]=16'he849;
aud[28510]=16'he85d;
aud[28511]=16'he871;
aud[28512]=16'he885;
aud[28513]=16'he899;
aud[28514]=16'he8ad;
aud[28515]=16'he8c0;
aud[28516]=16'he8d4;
aud[28517]=16'he8e8;
aud[28518]=16'he8fc;
aud[28519]=16'he910;
aud[28520]=16'he925;
aud[28521]=16'he939;
aud[28522]=16'he94d;
aud[28523]=16'he961;
aud[28524]=16'he975;
aud[28525]=16'he989;
aud[28526]=16'he99d;
aud[28527]=16'he9b1;
aud[28528]=16'he9c5;
aud[28529]=16'he9d9;
aud[28530]=16'he9ed;
aud[28531]=16'hea01;
aud[28532]=16'hea16;
aud[28533]=16'hea2a;
aud[28534]=16'hea3e;
aud[28535]=16'hea52;
aud[28536]=16'hea66;
aud[28537]=16'hea7a;
aud[28538]=16'hea8f;
aud[28539]=16'heaa3;
aud[28540]=16'heab7;
aud[28541]=16'heacb;
aud[28542]=16'heae0;
aud[28543]=16'heaf4;
aud[28544]=16'heb08;
aud[28545]=16'heb1c;
aud[28546]=16'heb31;
aud[28547]=16'heb45;
aud[28548]=16'heb59;
aud[28549]=16'heb6e;
aud[28550]=16'heb82;
aud[28551]=16'heb96;
aud[28552]=16'hebab;
aud[28553]=16'hebbf;
aud[28554]=16'hebd3;
aud[28555]=16'hebe8;
aud[28556]=16'hebfc;
aud[28557]=16'hec10;
aud[28558]=16'hec25;
aud[28559]=16'hec39;
aud[28560]=16'hec4d;
aud[28561]=16'hec62;
aud[28562]=16'hec76;
aud[28563]=16'hec8b;
aud[28564]=16'hec9f;
aud[28565]=16'hecb4;
aud[28566]=16'hecc8;
aud[28567]=16'hecdd;
aud[28568]=16'hecf1;
aud[28569]=16'hed05;
aud[28570]=16'hed1a;
aud[28571]=16'hed2e;
aud[28572]=16'hed43;
aud[28573]=16'hed57;
aud[28574]=16'hed6c;
aud[28575]=16'hed81;
aud[28576]=16'hed95;
aud[28577]=16'hedaa;
aud[28578]=16'hedbe;
aud[28579]=16'hedd3;
aud[28580]=16'hede7;
aud[28581]=16'hedfc;
aud[28582]=16'hee10;
aud[28583]=16'hee25;
aud[28584]=16'hee3a;
aud[28585]=16'hee4e;
aud[28586]=16'hee63;
aud[28587]=16'hee77;
aud[28588]=16'hee8c;
aud[28589]=16'heea1;
aud[28590]=16'heeb5;
aud[28591]=16'heeca;
aud[28592]=16'heedf;
aud[28593]=16'heef3;
aud[28594]=16'hef08;
aud[28595]=16'hef1d;
aud[28596]=16'hef31;
aud[28597]=16'hef46;
aud[28598]=16'hef5b;
aud[28599]=16'hef70;
aud[28600]=16'hef84;
aud[28601]=16'hef99;
aud[28602]=16'hefae;
aud[28603]=16'hefc2;
aud[28604]=16'hefd7;
aud[28605]=16'hefec;
aud[28606]=16'hf001;
aud[28607]=16'hf015;
aud[28608]=16'hf02a;
aud[28609]=16'hf03f;
aud[28610]=16'hf054;
aud[28611]=16'hf069;
aud[28612]=16'hf07d;
aud[28613]=16'hf092;
aud[28614]=16'hf0a7;
aud[28615]=16'hf0bc;
aud[28616]=16'hf0d1;
aud[28617]=16'hf0e6;
aud[28618]=16'hf0fa;
aud[28619]=16'hf10f;
aud[28620]=16'hf124;
aud[28621]=16'hf139;
aud[28622]=16'hf14e;
aud[28623]=16'hf163;
aud[28624]=16'hf178;
aud[28625]=16'hf18c;
aud[28626]=16'hf1a1;
aud[28627]=16'hf1b6;
aud[28628]=16'hf1cb;
aud[28629]=16'hf1e0;
aud[28630]=16'hf1f5;
aud[28631]=16'hf20a;
aud[28632]=16'hf21f;
aud[28633]=16'hf234;
aud[28634]=16'hf249;
aud[28635]=16'hf25e;
aud[28636]=16'hf273;
aud[28637]=16'hf288;
aud[28638]=16'hf29d;
aud[28639]=16'hf2b2;
aud[28640]=16'hf2c7;
aud[28641]=16'hf2dc;
aud[28642]=16'hf2f1;
aud[28643]=16'hf306;
aud[28644]=16'hf31b;
aud[28645]=16'hf330;
aud[28646]=16'hf345;
aud[28647]=16'hf35a;
aud[28648]=16'hf36f;
aud[28649]=16'hf384;
aud[28650]=16'hf399;
aud[28651]=16'hf3ae;
aud[28652]=16'hf3c3;
aud[28653]=16'hf3d8;
aud[28654]=16'hf3ed;
aud[28655]=16'hf402;
aud[28656]=16'hf417;
aud[28657]=16'hf42c;
aud[28658]=16'hf441;
aud[28659]=16'hf456;
aud[28660]=16'hf46b;
aud[28661]=16'hf480;
aud[28662]=16'hf496;
aud[28663]=16'hf4ab;
aud[28664]=16'hf4c0;
aud[28665]=16'hf4d5;
aud[28666]=16'hf4ea;
aud[28667]=16'hf4ff;
aud[28668]=16'hf514;
aud[28669]=16'hf529;
aud[28670]=16'hf53f;
aud[28671]=16'hf554;
aud[28672]=16'hf569;
aud[28673]=16'hf57e;
aud[28674]=16'hf593;
aud[28675]=16'hf5a8;
aud[28676]=16'hf5bd;
aud[28677]=16'hf5d3;
aud[28678]=16'hf5e8;
aud[28679]=16'hf5fd;
aud[28680]=16'hf612;
aud[28681]=16'hf627;
aud[28682]=16'hf63d;
aud[28683]=16'hf652;
aud[28684]=16'hf667;
aud[28685]=16'hf67c;
aud[28686]=16'hf691;
aud[28687]=16'hf6a7;
aud[28688]=16'hf6bc;
aud[28689]=16'hf6d1;
aud[28690]=16'hf6e6;
aud[28691]=16'hf6fb;
aud[28692]=16'hf711;
aud[28693]=16'hf726;
aud[28694]=16'hf73b;
aud[28695]=16'hf750;
aud[28696]=16'hf766;
aud[28697]=16'hf77b;
aud[28698]=16'hf790;
aud[28699]=16'hf7a5;
aud[28700]=16'hf7bb;
aud[28701]=16'hf7d0;
aud[28702]=16'hf7e5;
aud[28703]=16'hf7fb;
aud[28704]=16'hf810;
aud[28705]=16'hf825;
aud[28706]=16'hf83a;
aud[28707]=16'hf850;
aud[28708]=16'hf865;
aud[28709]=16'hf87a;
aud[28710]=16'hf890;
aud[28711]=16'hf8a5;
aud[28712]=16'hf8ba;
aud[28713]=16'hf8cf;
aud[28714]=16'hf8e5;
aud[28715]=16'hf8fa;
aud[28716]=16'hf90f;
aud[28717]=16'hf925;
aud[28718]=16'hf93a;
aud[28719]=16'hf94f;
aud[28720]=16'hf965;
aud[28721]=16'hf97a;
aud[28722]=16'hf98f;
aud[28723]=16'hf9a5;
aud[28724]=16'hf9ba;
aud[28725]=16'hf9cf;
aud[28726]=16'hf9e5;
aud[28727]=16'hf9fa;
aud[28728]=16'hfa0f;
aud[28729]=16'hfa25;
aud[28730]=16'hfa3a;
aud[28731]=16'hfa50;
aud[28732]=16'hfa65;
aud[28733]=16'hfa7a;
aud[28734]=16'hfa90;
aud[28735]=16'hfaa5;
aud[28736]=16'hfaba;
aud[28737]=16'hfad0;
aud[28738]=16'hfae5;
aud[28739]=16'hfafb;
aud[28740]=16'hfb10;
aud[28741]=16'hfb25;
aud[28742]=16'hfb3b;
aud[28743]=16'hfb50;
aud[28744]=16'hfb65;
aud[28745]=16'hfb7b;
aud[28746]=16'hfb90;
aud[28747]=16'hfba6;
aud[28748]=16'hfbbb;
aud[28749]=16'hfbd0;
aud[28750]=16'hfbe6;
aud[28751]=16'hfbfb;
aud[28752]=16'hfc11;
aud[28753]=16'hfc26;
aud[28754]=16'hfc3b;
aud[28755]=16'hfc51;
aud[28756]=16'hfc66;
aud[28757]=16'hfc7c;
aud[28758]=16'hfc91;
aud[28759]=16'hfca7;
aud[28760]=16'hfcbc;
aud[28761]=16'hfcd1;
aud[28762]=16'hfce7;
aud[28763]=16'hfcfc;
aud[28764]=16'hfd12;
aud[28765]=16'hfd27;
aud[28766]=16'hfd3c;
aud[28767]=16'hfd52;
aud[28768]=16'hfd67;
aud[28769]=16'hfd7d;
aud[28770]=16'hfd92;
aud[28771]=16'hfda8;
aud[28772]=16'hfdbd;
aud[28773]=16'hfdd2;
aud[28774]=16'hfde8;
aud[28775]=16'hfdfd;
aud[28776]=16'hfe13;
aud[28777]=16'hfe28;
aud[28778]=16'hfe3e;
aud[28779]=16'hfe53;
aud[28780]=16'hfe69;
aud[28781]=16'hfe7e;
aud[28782]=16'hfe93;
aud[28783]=16'hfea9;
aud[28784]=16'hfebe;
aud[28785]=16'hfed4;
aud[28786]=16'hfee9;
aud[28787]=16'hfeff;
aud[28788]=16'hff14;
aud[28789]=16'hff2a;
aud[28790]=16'hff3f;
aud[28791]=16'hff54;
aud[28792]=16'hff6a;
aud[28793]=16'hff7f;
aud[28794]=16'hff95;
aud[28795]=16'hffaa;
aud[28796]=16'hffc0;
aud[28797]=16'hffd5;
aud[28798]=16'hffeb;
aud[28799]=16'h0;
aud[28800]=16'h15;
aud[28801]=16'h2b;
aud[28802]=16'h40;
aud[28803]=16'h56;
aud[28804]=16'h6b;
aud[28805]=16'h81;
aud[28806]=16'h96;
aud[28807]=16'hac;
aud[28808]=16'hc1;
aud[28809]=16'hd6;
aud[28810]=16'hec;
aud[28811]=16'h101;
aud[28812]=16'h117;
aud[28813]=16'h12c;
aud[28814]=16'h142;
aud[28815]=16'h157;
aud[28816]=16'h16d;
aud[28817]=16'h182;
aud[28818]=16'h197;
aud[28819]=16'h1ad;
aud[28820]=16'h1c2;
aud[28821]=16'h1d8;
aud[28822]=16'h1ed;
aud[28823]=16'h203;
aud[28824]=16'h218;
aud[28825]=16'h22e;
aud[28826]=16'h243;
aud[28827]=16'h258;
aud[28828]=16'h26e;
aud[28829]=16'h283;
aud[28830]=16'h299;
aud[28831]=16'h2ae;
aud[28832]=16'h2c4;
aud[28833]=16'h2d9;
aud[28834]=16'h2ee;
aud[28835]=16'h304;
aud[28836]=16'h319;
aud[28837]=16'h32f;
aud[28838]=16'h344;
aud[28839]=16'h359;
aud[28840]=16'h36f;
aud[28841]=16'h384;
aud[28842]=16'h39a;
aud[28843]=16'h3af;
aud[28844]=16'h3c5;
aud[28845]=16'h3da;
aud[28846]=16'h3ef;
aud[28847]=16'h405;
aud[28848]=16'h41a;
aud[28849]=16'h430;
aud[28850]=16'h445;
aud[28851]=16'h45a;
aud[28852]=16'h470;
aud[28853]=16'h485;
aud[28854]=16'h49b;
aud[28855]=16'h4b0;
aud[28856]=16'h4c5;
aud[28857]=16'h4db;
aud[28858]=16'h4f0;
aud[28859]=16'h505;
aud[28860]=16'h51b;
aud[28861]=16'h530;
aud[28862]=16'h546;
aud[28863]=16'h55b;
aud[28864]=16'h570;
aud[28865]=16'h586;
aud[28866]=16'h59b;
aud[28867]=16'h5b0;
aud[28868]=16'h5c6;
aud[28869]=16'h5db;
aud[28870]=16'h5f1;
aud[28871]=16'h606;
aud[28872]=16'h61b;
aud[28873]=16'h631;
aud[28874]=16'h646;
aud[28875]=16'h65b;
aud[28876]=16'h671;
aud[28877]=16'h686;
aud[28878]=16'h69b;
aud[28879]=16'h6b1;
aud[28880]=16'h6c6;
aud[28881]=16'h6db;
aud[28882]=16'h6f1;
aud[28883]=16'h706;
aud[28884]=16'h71b;
aud[28885]=16'h731;
aud[28886]=16'h746;
aud[28887]=16'h75b;
aud[28888]=16'h770;
aud[28889]=16'h786;
aud[28890]=16'h79b;
aud[28891]=16'h7b0;
aud[28892]=16'h7c6;
aud[28893]=16'h7db;
aud[28894]=16'h7f0;
aud[28895]=16'h805;
aud[28896]=16'h81b;
aud[28897]=16'h830;
aud[28898]=16'h845;
aud[28899]=16'h85b;
aud[28900]=16'h870;
aud[28901]=16'h885;
aud[28902]=16'h89a;
aud[28903]=16'h8b0;
aud[28904]=16'h8c5;
aud[28905]=16'h8da;
aud[28906]=16'h8ef;
aud[28907]=16'h905;
aud[28908]=16'h91a;
aud[28909]=16'h92f;
aud[28910]=16'h944;
aud[28911]=16'h959;
aud[28912]=16'h96f;
aud[28913]=16'h984;
aud[28914]=16'h999;
aud[28915]=16'h9ae;
aud[28916]=16'h9c3;
aud[28917]=16'h9d9;
aud[28918]=16'h9ee;
aud[28919]=16'ha03;
aud[28920]=16'ha18;
aud[28921]=16'ha2d;
aud[28922]=16'ha43;
aud[28923]=16'ha58;
aud[28924]=16'ha6d;
aud[28925]=16'ha82;
aud[28926]=16'ha97;
aud[28927]=16'haac;
aud[28928]=16'hac1;
aud[28929]=16'had7;
aud[28930]=16'haec;
aud[28931]=16'hb01;
aud[28932]=16'hb16;
aud[28933]=16'hb2b;
aud[28934]=16'hb40;
aud[28935]=16'hb55;
aud[28936]=16'hb6a;
aud[28937]=16'hb80;
aud[28938]=16'hb95;
aud[28939]=16'hbaa;
aud[28940]=16'hbbf;
aud[28941]=16'hbd4;
aud[28942]=16'hbe9;
aud[28943]=16'hbfe;
aud[28944]=16'hc13;
aud[28945]=16'hc28;
aud[28946]=16'hc3d;
aud[28947]=16'hc52;
aud[28948]=16'hc67;
aud[28949]=16'hc7c;
aud[28950]=16'hc91;
aud[28951]=16'hca6;
aud[28952]=16'hcbb;
aud[28953]=16'hcd0;
aud[28954]=16'hce5;
aud[28955]=16'hcfa;
aud[28956]=16'hd0f;
aud[28957]=16'hd24;
aud[28958]=16'hd39;
aud[28959]=16'hd4e;
aud[28960]=16'hd63;
aud[28961]=16'hd78;
aud[28962]=16'hd8d;
aud[28963]=16'hda2;
aud[28964]=16'hdb7;
aud[28965]=16'hdcc;
aud[28966]=16'hde1;
aud[28967]=16'hdf6;
aud[28968]=16'he0b;
aud[28969]=16'he20;
aud[28970]=16'he35;
aud[28971]=16'he4a;
aud[28972]=16'he5f;
aud[28973]=16'he74;
aud[28974]=16'he88;
aud[28975]=16'he9d;
aud[28976]=16'heb2;
aud[28977]=16'hec7;
aud[28978]=16'hedc;
aud[28979]=16'hef1;
aud[28980]=16'hf06;
aud[28981]=16'hf1a;
aud[28982]=16'hf2f;
aud[28983]=16'hf44;
aud[28984]=16'hf59;
aud[28985]=16'hf6e;
aud[28986]=16'hf83;
aud[28987]=16'hf97;
aud[28988]=16'hfac;
aud[28989]=16'hfc1;
aud[28990]=16'hfd6;
aud[28991]=16'hfeb;
aud[28992]=16'hfff;
aud[28993]=16'h1014;
aud[28994]=16'h1029;
aud[28995]=16'h103e;
aud[28996]=16'h1052;
aud[28997]=16'h1067;
aud[28998]=16'h107c;
aud[28999]=16'h1090;
aud[29000]=16'h10a5;
aud[29001]=16'h10ba;
aud[29002]=16'h10cf;
aud[29003]=16'h10e3;
aud[29004]=16'h10f8;
aud[29005]=16'h110d;
aud[29006]=16'h1121;
aud[29007]=16'h1136;
aud[29008]=16'h114b;
aud[29009]=16'h115f;
aud[29010]=16'h1174;
aud[29011]=16'h1189;
aud[29012]=16'h119d;
aud[29013]=16'h11b2;
aud[29014]=16'h11c6;
aud[29015]=16'h11db;
aud[29016]=16'h11f0;
aud[29017]=16'h1204;
aud[29018]=16'h1219;
aud[29019]=16'h122d;
aud[29020]=16'h1242;
aud[29021]=16'h1256;
aud[29022]=16'h126b;
aud[29023]=16'h127f;
aud[29024]=16'h1294;
aud[29025]=16'h12a9;
aud[29026]=16'h12bd;
aud[29027]=16'h12d2;
aud[29028]=16'h12e6;
aud[29029]=16'h12fb;
aud[29030]=16'h130f;
aud[29031]=16'h1323;
aud[29032]=16'h1338;
aud[29033]=16'h134c;
aud[29034]=16'h1361;
aud[29035]=16'h1375;
aud[29036]=16'h138a;
aud[29037]=16'h139e;
aud[29038]=16'h13b3;
aud[29039]=16'h13c7;
aud[29040]=16'h13db;
aud[29041]=16'h13f0;
aud[29042]=16'h1404;
aud[29043]=16'h1418;
aud[29044]=16'h142d;
aud[29045]=16'h1441;
aud[29046]=16'h1455;
aud[29047]=16'h146a;
aud[29048]=16'h147e;
aud[29049]=16'h1492;
aud[29050]=16'h14a7;
aud[29051]=16'h14bb;
aud[29052]=16'h14cf;
aud[29053]=16'h14e4;
aud[29054]=16'h14f8;
aud[29055]=16'h150c;
aud[29056]=16'h1520;
aud[29057]=16'h1535;
aud[29058]=16'h1549;
aud[29059]=16'h155d;
aud[29060]=16'h1571;
aud[29061]=16'h1586;
aud[29062]=16'h159a;
aud[29063]=16'h15ae;
aud[29064]=16'h15c2;
aud[29065]=16'h15d6;
aud[29066]=16'h15ea;
aud[29067]=16'h15ff;
aud[29068]=16'h1613;
aud[29069]=16'h1627;
aud[29070]=16'h163b;
aud[29071]=16'h164f;
aud[29072]=16'h1663;
aud[29073]=16'h1677;
aud[29074]=16'h168b;
aud[29075]=16'h169f;
aud[29076]=16'h16b3;
aud[29077]=16'h16c7;
aud[29078]=16'h16db;
aud[29079]=16'h16f0;
aud[29080]=16'h1704;
aud[29081]=16'h1718;
aud[29082]=16'h172c;
aud[29083]=16'h1740;
aud[29084]=16'h1753;
aud[29085]=16'h1767;
aud[29086]=16'h177b;
aud[29087]=16'h178f;
aud[29088]=16'h17a3;
aud[29089]=16'h17b7;
aud[29090]=16'h17cb;
aud[29091]=16'h17df;
aud[29092]=16'h17f3;
aud[29093]=16'h1807;
aud[29094]=16'h181b;
aud[29095]=16'h182f;
aud[29096]=16'h1842;
aud[29097]=16'h1856;
aud[29098]=16'h186a;
aud[29099]=16'h187e;
aud[29100]=16'h1892;
aud[29101]=16'h18a5;
aud[29102]=16'h18b9;
aud[29103]=16'h18cd;
aud[29104]=16'h18e1;
aud[29105]=16'h18f5;
aud[29106]=16'h1908;
aud[29107]=16'h191c;
aud[29108]=16'h1930;
aud[29109]=16'h1943;
aud[29110]=16'h1957;
aud[29111]=16'h196b;
aud[29112]=16'h197f;
aud[29113]=16'h1992;
aud[29114]=16'h19a6;
aud[29115]=16'h19ba;
aud[29116]=16'h19cd;
aud[29117]=16'h19e1;
aud[29118]=16'h19f4;
aud[29119]=16'h1a08;
aud[29120]=16'h1a1c;
aud[29121]=16'h1a2f;
aud[29122]=16'h1a43;
aud[29123]=16'h1a56;
aud[29124]=16'h1a6a;
aud[29125]=16'h1a7d;
aud[29126]=16'h1a91;
aud[29127]=16'h1aa4;
aud[29128]=16'h1ab8;
aud[29129]=16'h1acb;
aud[29130]=16'h1adf;
aud[29131]=16'h1af2;
aud[29132]=16'h1b06;
aud[29133]=16'h1b19;
aud[29134]=16'h1b2d;
aud[29135]=16'h1b40;
aud[29136]=16'h1b53;
aud[29137]=16'h1b67;
aud[29138]=16'h1b7a;
aud[29139]=16'h1b8d;
aud[29140]=16'h1ba1;
aud[29141]=16'h1bb4;
aud[29142]=16'h1bc8;
aud[29143]=16'h1bdb;
aud[29144]=16'h1bee;
aud[29145]=16'h1c01;
aud[29146]=16'h1c15;
aud[29147]=16'h1c28;
aud[29148]=16'h1c3b;
aud[29149]=16'h1c4e;
aud[29150]=16'h1c62;
aud[29151]=16'h1c75;
aud[29152]=16'h1c88;
aud[29153]=16'h1c9b;
aud[29154]=16'h1cae;
aud[29155]=16'h1cc2;
aud[29156]=16'h1cd5;
aud[29157]=16'h1ce8;
aud[29158]=16'h1cfb;
aud[29159]=16'h1d0e;
aud[29160]=16'h1d21;
aud[29161]=16'h1d34;
aud[29162]=16'h1d47;
aud[29163]=16'h1d5b;
aud[29164]=16'h1d6e;
aud[29165]=16'h1d81;
aud[29166]=16'h1d94;
aud[29167]=16'h1da7;
aud[29168]=16'h1dba;
aud[29169]=16'h1dcd;
aud[29170]=16'h1de0;
aud[29171]=16'h1df3;
aud[29172]=16'h1e06;
aud[29173]=16'h1e18;
aud[29174]=16'h1e2b;
aud[29175]=16'h1e3e;
aud[29176]=16'h1e51;
aud[29177]=16'h1e64;
aud[29178]=16'h1e77;
aud[29179]=16'h1e8a;
aud[29180]=16'h1e9d;
aud[29181]=16'h1eaf;
aud[29182]=16'h1ec2;
aud[29183]=16'h1ed5;
aud[29184]=16'h1ee8;
aud[29185]=16'h1efb;
aud[29186]=16'h1f0d;
aud[29187]=16'h1f20;
aud[29188]=16'h1f33;
aud[29189]=16'h1f46;
aud[29190]=16'h1f58;
aud[29191]=16'h1f6b;
aud[29192]=16'h1f7e;
aud[29193]=16'h1f90;
aud[29194]=16'h1fa3;
aud[29195]=16'h1fb6;
aud[29196]=16'h1fc8;
aud[29197]=16'h1fdb;
aud[29198]=16'h1fed;
aud[29199]=16'h2000;
aud[29200]=16'h2013;
aud[29201]=16'h2025;
aud[29202]=16'h2038;
aud[29203]=16'h204a;
aud[29204]=16'h205d;
aud[29205]=16'h206f;
aud[29206]=16'h2082;
aud[29207]=16'h2094;
aud[29208]=16'h20a7;
aud[29209]=16'h20b9;
aud[29210]=16'h20cb;
aud[29211]=16'h20de;
aud[29212]=16'h20f0;
aud[29213]=16'h2103;
aud[29214]=16'h2115;
aud[29215]=16'h2127;
aud[29216]=16'h213a;
aud[29217]=16'h214c;
aud[29218]=16'h215e;
aud[29219]=16'h2171;
aud[29220]=16'h2183;
aud[29221]=16'h2195;
aud[29222]=16'h21a7;
aud[29223]=16'h21ba;
aud[29224]=16'h21cc;
aud[29225]=16'h21de;
aud[29226]=16'h21f0;
aud[29227]=16'h2202;
aud[29228]=16'h2215;
aud[29229]=16'h2227;
aud[29230]=16'h2239;
aud[29231]=16'h224b;
aud[29232]=16'h225d;
aud[29233]=16'h226f;
aud[29234]=16'h2281;
aud[29235]=16'h2293;
aud[29236]=16'h22a5;
aud[29237]=16'h22b7;
aud[29238]=16'h22c9;
aud[29239]=16'h22db;
aud[29240]=16'h22ed;
aud[29241]=16'h22ff;
aud[29242]=16'h2311;
aud[29243]=16'h2323;
aud[29244]=16'h2335;
aud[29245]=16'h2347;
aud[29246]=16'h2359;
aud[29247]=16'h236b;
aud[29248]=16'h237d;
aud[29249]=16'h238e;
aud[29250]=16'h23a0;
aud[29251]=16'h23b2;
aud[29252]=16'h23c4;
aud[29253]=16'h23d6;
aud[29254]=16'h23e7;
aud[29255]=16'h23f9;
aud[29256]=16'h240b;
aud[29257]=16'h241d;
aud[29258]=16'h242e;
aud[29259]=16'h2440;
aud[29260]=16'h2452;
aud[29261]=16'h2463;
aud[29262]=16'h2475;
aud[29263]=16'h2487;
aud[29264]=16'h2498;
aud[29265]=16'h24aa;
aud[29266]=16'h24bb;
aud[29267]=16'h24cd;
aud[29268]=16'h24de;
aud[29269]=16'h24f0;
aud[29270]=16'h2501;
aud[29271]=16'h2513;
aud[29272]=16'h2524;
aud[29273]=16'h2536;
aud[29274]=16'h2547;
aud[29275]=16'h2559;
aud[29276]=16'h256a;
aud[29277]=16'h257c;
aud[29278]=16'h258d;
aud[29279]=16'h259e;
aud[29280]=16'h25b0;
aud[29281]=16'h25c1;
aud[29282]=16'h25d2;
aud[29283]=16'h25e4;
aud[29284]=16'h25f5;
aud[29285]=16'h2606;
aud[29286]=16'h2617;
aud[29287]=16'h2629;
aud[29288]=16'h263a;
aud[29289]=16'h264b;
aud[29290]=16'h265c;
aud[29291]=16'h266d;
aud[29292]=16'h267e;
aud[29293]=16'h2690;
aud[29294]=16'h26a1;
aud[29295]=16'h26b2;
aud[29296]=16'h26c3;
aud[29297]=16'h26d4;
aud[29298]=16'h26e5;
aud[29299]=16'h26f6;
aud[29300]=16'h2707;
aud[29301]=16'h2718;
aud[29302]=16'h2729;
aud[29303]=16'h273a;
aud[29304]=16'h274b;
aud[29305]=16'h275c;
aud[29306]=16'h276d;
aud[29307]=16'h277e;
aud[29308]=16'h278e;
aud[29309]=16'h279f;
aud[29310]=16'h27b0;
aud[29311]=16'h27c1;
aud[29312]=16'h27d2;
aud[29313]=16'h27e2;
aud[29314]=16'h27f3;
aud[29315]=16'h2804;
aud[29316]=16'h2815;
aud[29317]=16'h2825;
aud[29318]=16'h2836;
aud[29319]=16'h2847;
aud[29320]=16'h2857;
aud[29321]=16'h2868;
aud[29322]=16'h2879;
aud[29323]=16'h2889;
aud[29324]=16'h289a;
aud[29325]=16'h28aa;
aud[29326]=16'h28bb;
aud[29327]=16'h28cc;
aud[29328]=16'h28dc;
aud[29329]=16'h28ed;
aud[29330]=16'h28fd;
aud[29331]=16'h290e;
aud[29332]=16'h291e;
aud[29333]=16'h292e;
aud[29334]=16'h293f;
aud[29335]=16'h294f;
aud[29336]=16'h2960;
aud[29337]=16'h2970;
aud[29338]=16'h2980;
aud[29339]=16'h2991;
aud[29340]=16'h29a1;
aud[29341]=16'h29b1;
aud[29342]=16'h29c1;
aud[29343]=16'h29d2;
aud[29344]=16'h29e2;
aud[29345]=16'h29f2;
aud[29346]=16'h2a02;
aud[29347]=16'h2a12;
aud[29348]=16'h2a23;
aud[29349]=16'h2a33;
aud[29350]=16'h2a43;
aud[29351]=16'h2a53;
aud[29352]=16'h2a63;
aud[29353]=16'h2a73;
aud[29354]=16'h2a83;
aud[29355]=16'h2a93;
aud[29356]=16'h2aa3;
aud[29357]=16'h2ab3;
aud[29358]=16'h2ac3;
aud[29359]=16'h2ad3;
aud[29360]=16'h2ae3;
aud[29361]=16'h2af3;
aud[29362]=16'h2b03;
aud[29363]=16'h2b13;
aud[29364]=16'h2b22;
aud[29365]=16'h2b32;
aud[29366]=16'h2b42;
aud[29367]=16'h2b52;
aud[29368]=16'h2b62;
aud[29369]=16'h2b71;
aud[29370]=16'h2b81;
aud[29371]=16'h2b91;
aud[29372]=16'h2ba1;
aud[29373]=16'h2bb0;
aud[29374]=16'h2bc0;
aud[29375]=16'h2bd0;
aud[29376]=16'h2bdf;
aud[29377]=16'h2bef;
aud[29378]=16'h2bfe;
aud[29379]=16'h2c0e;
aud[29380]=16'h2c1e;
aud[29381]=16'h2c2d;
aud[29382]=16'h2c3d;
aud[29383]=16'h2c4c;
aud[29384]=16'h2c5c;
aud[29385]=16'h2c6b;
aud[29386]=16'h2c7a;
aud[29387]=16'h2c8a;
aud[29388]=16'h2c99;
aud[29389]=16'h2ca9;
aud[29390]=16'h2cb8;
aud[29391]=16'h2cc7;
aud[29392]=16'h2cd7;
aud[29393]=16'h2ce6;
aud[29394]=16'h2cf5;
aud[29395]=16'h2d04;
aud[29396]=16'h2d14;
aud[29397]=16'h2d23;
aud[29398]=16'h2d32;
aud[29399]=16'h2d41;
aud[29400]=16'h2d50;
aud[29401]=16'h2d60;
aud[29402]=16'h2d6f;
aud[29403]=16'h2d7e;
aud[29404]=16'h2d8d;
aud[29405]=16'h2d9c;
aud[29406]=16'h2dab;
aud[29407]=16'h2dba;
aud[29408]=16'h2dc9;
aud[29409]=16'h2dd8;
aud[29410]=16'h2de7;
aud[29411]=16'h2df6;
aud[29412]=16'h2e05;
aud[29413]=16'h2e14;
aud[29414]=16'h2e22;
aud[29415]=16'h2e31;
aud[29416]=16'h2e40;
aud[29417]=16'h2e4f;
aud[29418]=16'h2e5e;
aud[29419]=16'h2e6d;
aud[29420]=16'h2e7b;
aud[29421]=16'h2e8a;
aud[29422]=16'h2e99;
aud[29423]=16'h2ea7;
aud[29424]=16'h2eb6;
aud[29425]=16'h2ec5;
aud[29426]=16'h2ed3;
aud[29427]=16'h2ee2;
aud[29428]=16'h2ef1;
aud[29429]=16'h2eff;
aud[29430]=16'h2f0e;
aud[29431]=16'h2f1c;
aud[29432]=16'h2f2b;
aud[29433]=16'h2f39;
aud[29434]=16'h2f48;
aud[29435]=16'h2f56;
aud[29436]=16'h2f65;
aud[29437]=16'h2f73;
aud[29438]=16'h2f81;
aud[29439]=16'h2f90;
aud[29440]=16'h2f9e;
aud[29441]=16'h2fac;
aud[29442]=16'h2fbb;
aud[29443]=16'h2fc9;
aud[29444]=16'h2fd7;
aud[29445]=16'h2fe5;
aud[29446]=16'h2ff4;
aud[29447]=16'h3002;
aud[29448]=16'h3010;
aud[29449]=16'h301e;
aud[29450]=16'h302c;
aud[29451]=16'h303a;
aud[29452]=16'h3048;
aud[29453]=16'h3057;
aud[29454]=16'h3065;
aud[29455]=16'h3073;
aud[29456]=16'h3081;
aud[29457]=16'h308f;
aud[29458]=16'h309d;
aud[29459]=16'h30aa;
aud[29460]=16'h30b8;
aud[29461]=16'h30c6;
aud[29462]=16'h30d4;
aud[29463]=16'h30e2;
aud[29464]=16'h30f0;
aud[29465]=16'h30fe;
aud[29466]=16'h310b;
aud[29467]=16'h3119;
aud[29468]=16'h3127;
aud[29469]=16'h3135;
aud[29470]=16'h3142;
aud[29471]=16'h3150;
aud[29472]=16'h315e;
aud[29473]=16'h316b;
aud[29474]=16'h3179;
aud[29475]=16'h3187;
aud[29476]=16'h3194;
aud[29477]=16'h31a2;
aud[29478]=16'h31af;
aud[29479]=16'h31bd;
aud[29480]=16'h31ca;
aud[29481]=16'h31d8;
aud[29482]=16'h31e5;
aud[29483]=16'h31f3;
aud[29484]=16'h3200;
aud[29485]=16'h320d;
aud[29486]=16'h321b;
aud[29487]=16'h3228;
aud[29488]=16'h3235;
aud[29489]=16'h3243;
aud[29490]=16'h3250;
aud[29491]=16'h325d;
aud[29492]=16'h326a;
aud[29493]=16'h3278;
aud[29494]=16'h3285;
aud[29495]=16'h3292;
aud[29496]=16'h329f;
aud[29497]=16'h32ac;
aud[29498]=16'h32b9;
aud[29499]=16'h32c6;
aud[29500]=16'h32d3;
aud[29501]=16'h32e0;
aud[29502]=16'h32ed;
aud[29503]=16'h32fa;
aud[29504]=16'h3307;
aud[29505]=16'h3314;
aud[29506]=16'h3321;
aud[29507]=16'h332e;
aud[29508]=16'h333b;
aud[29509]=16'h3348;
aud[29510]=16'h3355;
aud[29511]=16'h3361;
aud[29512]=16'h336e;
aud[29513]=16'h337b;
aud[29514]=16'h3388;
aud[29515]=16'h3394;
aud[29516]=16'h33a1;
aud[29517]=16'h33ae;
aud[29518]=16'h33ba;
aud[29519]=16'h33c7;
aud[29520]=16'h33d4;
aud[29521]=16'h33e0;
aud[29522]=16'h33ed;
aud[29523]=16'h33f9;
aud[29524]=16'h3406;
aud[29525]=16'h3412;
aud[29526]=16'h341f;
aud[29527]=16'h342b;
aud[29528]=16'h3437;
aud[29529]=16'h3444;
aud[29530]=16'h3450;
aud[29531]=16'h345d;
aud[29532]=16'h3469;
aud[29533]=16'h3475;
aud[29534]=16'h3481;
aud[29535]=16'h348e;
aud[29536]=16'h349a;
aud[29537]=16'h34a6;
aud[29538]=16'h34b2;
aud[29539]=16'h34be;
aud[29540]=16'h34cb;
aud[29541]=16'h34d7;
aud[29542]=16'h34e3;
aud[29543]=16'h34ef;
aud[29544]=16'h34fb;
aud[29545]=16'h3507;
aud[29546]=16'h3513;
aud[29547]=16'h351f;
aud[29548]=16'h352b;
aud[29549]=16'h3537;
aud[29550]=16'h3543;
aud[29551]=16'h354f;
aud[29552]=16'h355a;
aud[29553]=16'h3566;
aud[29554]=16'h3572;
aud[29555]=16'h357e;
aud[29556]=16'h358a;
aud[29557]=16'h3595;
aud[29558]=16'h35a1;
aud[29559]=16'h35ad;
aud[29560]=16'h35b8;
aud[29561]=16'h35c4;
aud[29562]=16'h35d0;
aud[29563]=16'h35db;
aud[29564]=16'h35e7;
aud[29565]=16'h35f2;
aud[29566]=16'h35fe;
aud[29567]=16'h3609;
aud[29568]=16'h3615;
aud[29569]=16'h3620;
aud[29570]=16'h362c;
aud[29571]=16'h3637;
aud[29572]=16'h3643;
aud[29573]=16'h364e;
aud[29574]=16'h3659;
aud[29575]=16'h3665;
aud[29576]=16'h3670;
aud[29577]=16'h367b;
aud[29578]=16'h3686;
aud[29579]=16'h3692;
aud[29580]=16'h369d;
aud[29581]=16'h36a8;
aud[29582]=16'h36b3;
aud[29583]=16'h36be;
aud[29584]=16'h36c9;
aud[29585]=16'h36d4;
aud[29586]=16'h36e0;
aud[29587]=16'h36eb;
aud[29588]=16'h36f6;
aud[29589]=16'h3701;
aud[29590]=16'h370b;
aud[29591]=16'h3716;
aud[29592]=16'h3721;
aud[29593]=16'h372c;
aud[29594]=16'h3737;
aud[29595]=16'h3742;
aud[29596]=16'h374d;
aud[29597]=16'h3757;
aud[29598]=16'h3762;
aud[29599]=16'h376d;
aud[29600]=16'h3778;
aud[29601]=16'h3782;
aud[29602]=16'h378d;
aud[29603]=16'h3798;
aud[29604]=16'h37a2;
aud[29605]=16'h37ad;
aud[29606]=16'h37b7;
aud[29607]=16'h37c2;
aud[29608]=16'h37cc;
aud[29609]=16'h37d7;
aud[29610]=16'h37e1;
aud[29611]=16'h37ec;
aud[29612]=16'h37f6;
aud[29613]=16'h3801;
aud[29614]=16'h380b;
aud[29615]=16'h3815;
aud[29616]=16'h3820;
aud[29617]=16'h382a;
aud[29618]=16'h3834;
aud[29619]=16'h383f;
aud[29620]=16'h3849;
aud[29621]=16'h3853;
aud[29622]=16'h385d;
aud[29623]=16'h3867;
aud[29624]=16'h3871;
aud[29625]=16'h387b;
aud[29626]=16'h3886;
aud[29627]=16'h3890;
aud[29628]=16'h389a;
aud[29629]=16'h38a4;
aud[29630]=16'h38ae;
aud[29631]=16'h38b8;
aud[29632]=16'h38c1;
aud[29633]=16'h38cb;
aud[29634]=16'h38d5;
aud[29635]=16'h38df;
aud[29636]=16'h38e9;
aud[29637]=16'h38f3;
aud[29638]=16'h38fd;
aud[29639]=16'h3906;
aud[29640]=16'h3910;
aud[29641]=16'h391a;
aud[29642]=16'h3923;
aud[29643]=16'h392d;
aud[29644]=16'h3937;
aud[29645]=16'h3940;
aud[29646]=16'h394a;
aud[29647]=16'h3953;
aud[29648]=16'h395d;
aud[29649]=16'h3966;
aud[29650]=16'h3970;
aud[29651]=16'h3979;
aud[29652]=16'h3983;
aud[29653]=16'h398c;
aud[29654]=16'h3995;
aud[29655]=16'h399f;
aud[29656]=16'h39a8;
aud[29657]=16'h39b1;
aud[29658]=16'h39bb;
aud[29659]=16'h39c4;
aud[29660]=16'h39cd;
aud[29661]=16'h39d6;
aud[29662]=16'h39e0;
aud[29663]=16'h39e9;
aud[29664]=16'h39f2;
aud[29665]=16'h39fb;
aud[29666]=16'h3a04;
aud[29667]=16'h3a0d;
aud[29668]=16'h3a16;
aud[29669]=16'h3a1f;
aud[29670]=16'h3a28;
aud[29671]=16'h3a31;
aud[29672]=16'h3a3a;
aud[29673]=16'h3a43;
aud[29674]=16'h3a4c;
aud[29675]=16'h3a54;
aud[29676]=16'h3a5d;
aud[29677]=16'h3a66;
aud[29678]=16'h3a6f;
aud[29679]=16'h3a78;
aud[29680]=16'h3a80;
aud[29681]=16'h3a89;
aud[29682]=16'h3a92;
aud[29683]=16'h3a9a;
aud[29684]=16'h3aa3;
aud[29685]=16'h3aab;
aud[29686]=16'h3ab4;
aud[29687]=16'h3abc;
aud[29688]=16'h3ac5;
aud[29689]=16'h3acd;
aud[29690]=16'h3ad6;
aud[29691]=16'h3ade;
aud[29692]=16'h3ae7;
aud[29693]=16'h3aef;
aud[29694]=16'h3af7;
aud[29695]=16'h3b00;
aud[29696]=16'h3b08;
aud[29697]=16'h3b10;
aud[29698]=16'h3b19;
aud[29699]=16'h3b21;
aud[29700]=16'h3b29;
aud[29701]=16'h3b31;
aud[29702]=16'h3b39;
aud[29703]=16'h3b41;
aud[29704]=16'h3b4a;
aud[29705]=16'h3b52;
aud[29706]=16'h3b5a;
aud[29707]=16'h3b62;
aud[29708]=16'h3b6a;
aud[29709]=16'h3b72;
aud[29710]=16'h3b7a;
aud[29711]=16'h3b81;
aud[29712]=16'h3b89;
aud[29713]=16'h3b91;
aud[29714]=16'h3b99;
aud[29715]=16'h3ba1;
aud[29716]=16'h3ba9;
aud[29717]=16'h3bb0;
aud[29718]=16'h3bb8;
aud[29719]=16'h3bc0;
aud[29720]=16'h3bc7;
aud[29721]=16'h3bcf;
aud[29722]=16'h3bd7;
aud[29723]=16'h3bde;
aud[29724]=16'h3be6;
aud[29725]=16'h3bed;
aud[29726]=16'h3bf5;
aud[29727]=16'h3bfc;
aud[29728]=16'h3c04;
aud[29729]=16'h3c0b;
aud[29730]=16'h3c13;
aud[29731]=16'h3c1a;
aud[29732]=16'h3c21;
aud[29733]=16'h3c29;
aud[29734]=16'h3c30;
aud[29735]=16'h3c37;
aud[29736]=16'h3c3f;
aud[29737]=16'h3c46;
aud[29738]=16'h3c4d;
aud[29739]=16'h3c54;
aud[29740]=16'h3c5b;
aud[29741]=16'h3c63;
aud[29742]=16'h3c6a;
aud[29743]=16'h3c71;
aud[29744]=16'h3c78;
aud[29745]=16'h3c7f;
aud[29746]=16'h3c86;
aud[29747]=16'h3c8d;
aud[29748]=16'h3c94;
aud[29749]=16'h3c9b;
aud[29750]=16'h3ca1;
aud[29751]=16'h3ca8;
aud[29752]=16'h3caf;
aud[29753]=16'h3cb6;
aud[29754]=16'h3cbd;
aud[29755]=16'h3cc3;
aud[29756]=16'h3cca;
aud[29757]=16'h3cd1;
aud[29758]=16'h3cd7;
aud[29759]=16'h3cde;
aud[29760]=16'h3ce5;
aud[29761]=16'h3ceb;
aud[29762]=16'h3cf2;
aud[29763]=16'h3cf8;
aud[29764]=16'h3cff;
aud[29765]=16'h3d05;
aud[29766]=16'h3d0c;
aud[29767]=16'h3d12;
aud[29768]=16'h3d19;
aud[29769]=16'h3d1f;
aud[29770]=16'h3d25;
aud[29771]=16'h3d2c;
aud[29772]=16'h3d32;
aud[29773]=16'h3d38;
aud[29774]=16'h3d3f;
aud[29775]=16'h3d45;
aud[29776]=16'h3d4b;
aud[29777]=16'h3d51;
aud[29778]=16'h3d57;
aud[29779]=16'h3d5d;
aud[29780]=16'h3d63;
aud[29781]=16'h3d69;
aud[29782]=16'h3d6f;
aud[29783]=16'h3d75;
aud[29784]=16'h3d7b;
aud[29785]=16'h3d81;
aud[29786]=16'h3d87;
aud[29787]=16'h3d8d;
aud[29788]=16'h3d93;
aud[29789]=16'h3d99;
aud[29790]=16'h3d9f;
aud[29791]=16'h3da4;
aud[29792]=16'h3daa;
aud[29793]=16'h3db0;
aud[29794]=16'h3db6;
aud[29795]=16'h3dbb;
aud[29796]=16'h3dc1;
aud[29797]=16'h3dc7;
aud[29798]=16'h3dcc;
aud[29799]=16'h3dd2;
aud[29800]=16'h3dd7;
aud[29801]=16'h3ddd;
aud[29802]=16'h3de2;
aud[29803]=16'h3de8;
aud[29804]=16'h3ded;
aud[29805]=16'h3df3;
aud[29806]=16'h3df8;
aud[29807]=16'h3dfd;
aud[29808]=16'h3e03;
aud[29809]=16'h3e08;
aud[29810]=16'h3e0d;
aud[29811]=16'h3e12;
aud[29812]=16'h3e18;
aud[29813]=16'h3e1d;
aud[29814]=16'h3e22;
aud[29815]=16'h3e27;
aud[29816]=16'h3e2c;
aud[29817]=16'h3e31;
aud[29818]=16'h3e36;
aud[29819]=16'h3e3b;
aud[29820]=16'h3e40;
aud[29821]=16'h3e45;
aud[29822]=16'h3e4a;
aud[29823]=16'h3e4f;
aud[29824]=16'h3e54;
aud[29825]=16'h3e59;
aud[29826]=16'h3e5e;
aud[29827]=16'h3e62;
aud[29828]=16'h3e67;
aud[29829]=16'h3e6c;
aud[29830]=16'h3e71;
aud[29831]=16'h3e75;
aud[29832]=16'h3e7a;
aud[29833]=16'h3e7f;
aud[29834]=16'h3e83;
aud[29835]=16'h3e88;
aud[29836]=16'h3e8c;
aud[29837]=16'h3e91;
aud[29838]=16'h3e95;
aud[29839]=16'h3e9a;
aud[29840]=16'h3e9e;
aud[29841]=16'h3ea3;
aud[29842]=16'h3ea7;
aud[29843]=16'h3eac;
aud[29844]=16'h3eb0;
aud[29845]=16'h3eb4;
aud[29846]=16'h3eb9;
aud[29847]=16'h3ebd;
aud[29848]=16'h3ec1;
aud[29849]=16'h3ec5;
aud[29850]=16'h3ec9;
aud[29851]=16'h3ecd;
aud[29852]=16'h3ed2;
aud[29853]=16'h3ed6;
aud[29854]=16'h3eda;
aud[29855]=16'h3ede;
aud[29856]=16'h3ee2;
aud[29857]=16'h3ee6;
aud[29858]=16'h3eea;
aud[29859]=16'h3eee;
aud[29860]=16'h3ef2;
aud[29861]=16'h3ef5;
aud[29862]=16'h3ef9;
aud[29863]=16'h3efd;
aud[29864]=16'h3f01;
aud[29865]=16'h3f05;
aud[29866]=16'h3f08;
aud[29867]=16'h3f0c;
aud[29868]=16'h3f10;
aud[29869]=16'h3f13;
aud[29870]=16'h3f17;
aud[29871]=16'h3f1b;
aud[29872]=16'h3f1e;
aud[29873]=16'h3f22;
aud[29874]=16'h3f25;
aud[29875]=16'h3f29;
aud[29876]=16'h3f2c;
aud[29877]=16'h3f30;
aud[29878]=16'h3f33;
aud[29879]=16'h3f36;
aud[29880]=16'h3f3a;
aud[29881]=16'h3f3d;
aud[29882]=16'h3f40;
aud[29883]=16'h3f43;
aud[29884]=16'h3f47;
aud[29885]=16'h3f4a;
aud[29886]=16'h3f4d;
aud[29887]=16'h3f50;
aud[29888]=16'h3f53;
aud[29889]=16'h3f56;
aud[29890]=16'h3f5a;
aud[29891]=16'h3f5d;
aud[29892]=16'h3f60;
aud[29893]=16'h3f63;
aud[29894]=16'h3f65;
aud[29895]=16'h3f68;
aud[29896]=16'h3f6b;
aud[29897]=16'h3f6e;
aud[29898]=16'h3f71;
aud[29899]=16'h3f74;
aud[29900]=16'h3f77;
aud[29901]=16'h3f79;
aud[29902]=16'h3f7c;
aud[29903]=16'h3f7f;
aud[29904]=16'h3f81;
aud[29905]=16'h3f84;
aud[29906]=16'h3f87;
aud[29907]=16'h3f89;
aud[29908]=16'h3f8c;
aud[29909]=16'h3f8e;
aud[29910]=16'h3f91;
aud[29911]=16'h3f93;
aud[29912]=16'h3f96;
aud[29913]=16'h3f98;
aud[29914]=16'h3f9b;
aud[29915]=16'h3f9d;
aud[29916]=16'h3f9f;
aud[29917]=16'h3fa2;
aud[29918]=16'h3fa4;
aud[29919]=16'h3fa6;
aud[29920]=16'h3fa8;
aud[29921]=16'h3fab;
aud[29922]=16'h3fad;
aud[29923]=16'h3faf;
aud[29924]=16'h3fb1;
aud[29925]=16'h3fb3;
aud[29926]=16'h3fb5;
aud[29927]=16'h3fb7;
aud[29928]=16'h3fb9;
aud[29929]=16'h3fbb;
aud[29930]=16'h3fbd;
aud[29931]=16'h3fbf;
aud[29932]=16'h3fc1;
aud[29933]=16'h3fc3;
aud[29934]=16'h3fc5;
aud[29935]=16'h3fc7;
aud[29936]=16'h3fc8;
aud[29937]=16'h3fca;
aud[29938]=16'h3fcc;
aud[29939]=16'h3fcd;
aud[29940]=16'h3fcf;
aud[29941]=16'h3fd1;
aud[29942]=16'h3fd2;
aud[29943]=16'h3fd4;
aud[29944]=16'h3fd6;
aud[29945]=16'h3fd7;
aud[29946]=16'h3fd9;
aud[29947]=16'h3fda;
aud[29948]=16'h3fdc;
aud[29949]=16'h3fdd;
aud[29950]=16'h3fde;
aud[29951]=16'h3fe0;
aud[29952]=16'h3fe1;
aud[29953]=16'h3fe2;
aud[29954]=16'h3fe4;
aud[29955]=16'h3fe5;
aud[29956]=16'h3fe6;
aud[29957]=16'h3fe7;
aud[29958]=16'h3fe8;
aud[29959]=16'h3fea;
aud[29960]=16'h3feb;
aud[29961]=16'h3fec;
aud[29962]=16'h3fed;
aud[29963]=16'h3fee;
aud[29964]=16'h3fef;
aud[29965]=16'h3ff0;
aud[29966]=16'h3ff1;
aud[29967]=16'h3ff2;
aud[29968]=16'h3ff3;
aud[29969]=16'h3ff3;
aud[29970]=16'h3ff4;
aud[29971]=16'h3ff5;
aud[29972]=16'h3ff6;
aud[29973]=16'h3ff7;
aud[29974]=16'h3ff7;
aud[29975]=16'h3ff8;
aud[29976]=16'h3ff9;
aud[29977]=16'h3ff9;
aud[29978]=16'h3ffa;
aud[29979]=16'h3ffa;
aud[29980]=16'h3ffb;
aud[29981]=16'h3ffb;
aud[29982]=16'h3ffc;
aud[29983]=16'h3ffc;
aud[29984]=16'h3ffd;
aud[29985]=16'h3ffd;
aud[29986]=16'h3ffe;
aud[29987]=16'h3ffe;
aud[29988]=16'h3ffe;
aud[29989]=16'h3fff;
aud[29990]=16'h3fff;
aud[29991]=16'h3fff;
aud[29992]=16'h3fff;
aud[29993]=16'h3fff;
aud[29994]=16'h4000;
aud[29995]=16'h4000;
aud[29996]=16'h4000;
aud[29997]=16'h4000;
aud[29998]=16'h4000;
aud[29999]=16'h4000;
aud[30000]=16'h4000;
aud[30001]=16'h4000;
aud[30002]=16'h4000;
aud[30003]=16'h4000;
aud[30004]=16'h4000;
aud[30005]=16'h3fff;
aud[30006]=16'h3fff;
aud[30007]=16'h3fff;
aud[30008]=16'h3fff;
aud[30009]=16'h3fff;
aud[30010]=16'h3ffe;
aud[30011]=16'h3ffe;
aud[30012]=16'h3ffe;
aud[30013]=16'h3ffd;
aud[30014]=16'h3ffd;
aud[30015]=16'h3ffc;
aud[30016]=16'h3ffc;
aud[30017]=16'h3ffb;
aud[30018]=16'h3ffb;
aud[30019]=16'h3ffa;
aud[30020]=16'h3ffa;
aud[30021]=16'h3ff9;
aud[30022]=16'h3ff9;
aud[30023]=16'h3ff8;
aud[30024]=16'h3ff7;
aud[30025]=16'h3ff7;
aud[30026]=16'h3ff6;
aud[30027]=16'h3ff5;
aud[30028]=16'h3ff4;
aud[30029]=16'h3ff3;
aud[30030]=16'h3ff3;
aud[30031]=16'h3ff2;
aud[30032]=16'h3ff1;
aud[30033]=16'h3ff0;
aud[30034]=16'h3fef;
aud[30035]=16'h3fee;
aud[30036]=16'h3fed;
aud[30037]=16'h3fec;
aud[30038]=16'h3feb;
aud[30039]=16'h3fea;
aud[30040]=16'h3fe8;
aud[30041]=16'h3fe7;
aud[30042]=16'h3fe6;
aud[30043]=16'h3fe5;
aud[30044]=16'h3fe4;
aud[30045]=16'h3fe2;
aud[30046]=16'h3fe1;
aud[30047]=16'h3fe0;
aud[30048]=16'h3fde;
aud[30049]=16'h3fdd;
aud[30050]=16'h3fdc;
aud[30051]=16'h3fda;
aud[30052]=16'h3fd9;
aud[30053]=16'h3fd7;
aud[30054]=16'h3fd6;
aud[30055]=16'h3fd4;
aud[30056]=16'h3fd2;
aud[30057]=16'h3fd1;
aud[30058]=16'h3fcf;
aud[30059]=16'h3fcd;
aud[30060]=16'h3fcc;
aud[30061]=16'h3fca;
aud[30062]=16'h3fc8;
aud[30063]=16'h3fc7;
aud[30064]=16'h3fc5;
aud[30065]=16'h3fc3;
aud[30066]=16'h3fc1;
aud[30067]=16'h3fbf;
aud[30068]=16'h3fbd;
aud[30069]=16'h3fbb;
aud[30070]=16'h3fb9;
aud[30071]=16'h3fb7;
aud[30072]=16'h3fb5;
aud[30073]=16'h3fb3;
aud[30074]=16'h3fb1;
aud[30075]=16'h3faf;
aud[30076]=16'h3fad;
aud[30077]=16'h3fab;
aud[30078]=16'h3fa8;
aud[30079]=16'h3fa6;
aud[30080]=16'h3fa4;
aud[30081]=16'h3fa2;
aud[30082]=16'h3f9f;
aud[30083]=16'h3f9d;
aud[30084]=16'h3f9b;
aud[30085]=16'h3f98;
aud[30086]=16'h3f96;
aud[30087]=16'h3f93;
aud[30088]=16'h3f91;
aud[30089]=16'h3f8e;
aud[30090]=16'h3f8c;
aud[30091]=16'h3f89;
aud[30092]=16'h3f87;
aud[30093]=16'h3f84;
aud[30094]=16'h3f81;
aud[30095]=16'h3f7f;
aud[30096]=16'h3f7c;
aud[30097]=16'h3f79;
aud[30098]=16'h3f77;
aud[30099]=16'h3f74;
aud[30100]=16'h3f71;
aud[30101]=16'h3f6e;
aud[30102]=16'h3f6b;
aud[30103]=16'h3f68;
aud[30104]=16'h3f65;
aud[30105]=16'h3f63;
aud[30106]=16'h3f60;
aud[30107]=16'h3f5d;
aud[30108]=16'h3f5a;
aud[30109]=16'h3f56;
aud[30110]=16'h3f53;
aud[30111]=16'h3f50;
aud[30112]=16'h3f4d;
aud[30113]=16'h3f4a;
aud[30114]=16'h3f47;
aud[30115]=16'h3f43;
aud[30116]=16'h3f40;
aud[30117]=16'h3f3d;
aud[30118]=16'h3f3a;
aud[30119]=16'h3f36;
aud[30120]=16'h3f33;
aud[30121]=16'h3f30;
aud[30122]=16'h3f2c;
aud[30123]=16'h3f29;
aud[30124]=16'h3f25;
aud[30125]=16'h3f22;
aud[30126]=16'h3f1e;
aud[30127]=16'h3f1b;
aud[30128]=16'h3f17;
aud[30129]=16'h3f13;
aud[30130]=16'h3f10;
aud[30131]=16'h3f0c;
aud[30132]=16'h3f08;
aud[30133]=16'h3f05;
aud[30134]=16'h3f01;
aud[30135]=16'h3efd;
aud[30136]=16'h3ef9;
aud[30137]=16'h3ef5;
aud[30138]=16'h3ef2;
aud[30139]=16'h3eee;
aud[30140]=16'h3eea;
aud[30141]=16'h3ee6;
aud[30142]=16'h3ee2;
aud[30143]=16'h3ede;
aud[30144]=16'h3eda;
aud[30145]=16'h3ed6;
aud[30146]=16'h3ed2;
aud[30147]=16'h3ecd;
aud[30148]=16'h3ec9;
aud[30149]=16'h3ec5;
aud[30150]=16'h3ec1;
aud[30151]=16'h3ebd;
aud[30152]=16'h3eb9;
aud[30153]=16'h3eb4;
aud[30154]=16'h3eb0;
aud[30155]=16'h3eac;
aud[30156]=16'h3ea7;
aud[30157]=16'h3ea3;
aud[30158]=16'h3e9e;
aud[30159]=16'h3e9a;
aud[30160]=16'h3e95;
aud[30161]=16'h3e91;
aud[30162]=16'h3e8c;
aud[30163]=16'h3e88;
aud[30164]=16'h3e83;
aud[30165]=16'h3e7f;
aud[30166]=16'h3e7a;
aud[30167]=16'h3e75;
aud[30168]=16'h3e71;
aud[30169]=16'h3e6c;
aud[30170]=16'h3e67;
aud[30171]=16'h3e62;
aud[30172]=16'h3e5e;
aud[30173]=16'h3e59;
aud[30174]=16'h3e54;
aud[30175]=16'h3e4f;
aud[30176]=16'h3e4a;
aud[30177]=16'h3e45;
aud[30178]=16'h3e40;
aud[30179]=16'h3e3b;
aud[30180]=16'h3e36;
aud[30181]=16'h3e31;
aud[30182]=16'h3e2c;
aud[30183]=16'h3e27;
aud[30184]=16'h3e22;
aud[30185]=16'h3e1d;
aud[30186]=16'h3e18;
aud[30187]=16'h3e12;
aud[30188]=16'h3e0d;
aud[30189]=16'h3e08;
aud[30190]=16'h3e03;
aud[30191]=16'h3dfd;
aud[30192]=16'h3df8;
aud[30193]=16'h3df3;
aud[30194]=16'h3ded;
aud[30195]=16'h3de8;
aud[30196]=16'h3de2;
aud[30197]=16'h3ddd;
aud[30198]=16'h3dd7;
aud[30199]=16'h3dd2;
aud[30200]=16'h3dcc;
aud[30201]=16'h3dc7;
aud[30202]=16'h3dc1;
aud[30203]=16'h3dbb;
aud[30204]=16'h3db6;
aud[30205]=16'h3db0;
aud[30206]=16'h3daa;
aud[30207]=16'h3da4;
aud[30208]=16'h3d9f;
aud[30209]=16'h3d99;
aud[30210]=16'h3d93;
aud[30211]=16'h3d8d;
aud[30212]=16'h3d87;
aud[30213]=16'h3d81;
aud[30214]=16'h3d7b;
aud[30215]=16'h3d75;
aud[30216]=16'h3d6f;
aud[30217]=16'h3d69;
aud[30218]=16'h3d63;
aud[30219]=16'h3d5d;
aud[30220]=16'h3d57;
aud[30221]=16'h3d51;
aud[30222]=16'h3d4b;
aud[30223]=16'h3d45;
aud[30224]=16'h3d3f;
aud[30225]=16'h3d38;
aud[30226]=16'h3d32;
aud[30227]=16'h3d2c;
aud[30228]=16'h3d25;
aud[30229]=16'h3d1f;
aud[30230]=16'h3d19;
aud[30231]=16'h3d12;
aud[30232]=16'h3d0c;
aud[30233]=16'h3d05;
aud[30234]=16'h3cff;
aud[30235]=16'h3cf8;
aud[30236]=16'h3cf2;
aud[30237]=16'h3ceb;
aud[30238]=16'h3ce5;
aud[30239]=16'h3cde;
aud[30240]=16'h3cd7;
aud[30241]=16'h3cd1;
aud[30242]=16'h3cca;
aud[30243]=16'h3cc3;
aud[30244]=16'h3cbd;
aud[30245]=16'h3cb6;
aud[30246]=16'h3caf;
aud[30247]=16'h3ca8;
aud[30248]=16'h3ca1;
aud[30249]=16'h3c9b;
aud[30250]=16'h3c94;
aud[30251]=16'h3c8d;
aud[30252]=16'h3c86;
aud[30253]=16'h3c7f;
aud[30254]=16'h3c78;
aud[30255]=16'h3c71;
aud[30256]=16'h3c6a;
aud[30257]=16'h3c63;
aud[30258]=16'h3c5b;
aud[30259]=16'h3c54;
aud[30260]=16'h3c4d;
aud[30261]=16'h3c46;
aud[30262]=16'h3c3f;
aud[30263]=16'h3c37;
aud[30264]=16'h3c30;
aud[30265]=16'h3c29;
aud[30266]=16'h3c21;
aud[30267]=16'h3c1a;
aud[30268]=16'h3c13;
aud[30269]=16'h3c0b;
aud[30270]=16'h3c04;
aud[30271]=16'h3bfc;
aud[30272]=16'h3bf5;
aud[30273]=16'h3bed;
aud[30274]=16'h3be6;
aud[30275]=16'h3bde;
aud[30276]=16'h3bd7;
aud[30277]=16'h3bcf;
aud[30278]=16'h3bc7;
aud[30279]=16'h3bc0;
aud[30280]=16'h3bb8;
aud[30281]=16'h3bb0;
aud[30282]=16'h3ba9;
aud[30283]=16'h3ba1;
aud[30284]=16'h3b99;
aud[30285]=16'h3b91;
aud[30286]=16'h3b89;
aud[30287]=16'h3b81;
aud[30288]=16'h3b7a;
aud[30289]=16'h3b72;
aud[30290]=16'h3b6a;
aud[30291]=16'h3b62;
aud[30292]=16'h3b5a;
aud[30293]=16'h3b52;
aud[30294]=16'h3b4a;
aud[30295]=16'h3b41;
aud[30296]=16'h3b39;
aud[30297]=16'h3b31;
aud[30298]=16'h3b29;
aud[30299]=16'h3b21;
aud[30300]=16'h3b19;
aud[30301]=16'h3b10;
aud[30302]=16'h3b08;
aud[30303]=16'h3b00;
aud[30304]=16'h3af7;
aud[30305]=16'h3aef;
aud[30306]=16'h3ae7;
aud[30307]=16'h3ade;
aud[30308]=16'h3ad6;
aud[30309]=16'h3acd;
aud[30310]=16'h3ac5;
aud[30311]=16'h3abc;
aud[30312]=16'h3ab4;
aud[30313]=16'h3aab;
aud[30314]=16'h3aa3;
aud[30315]=16'h3a9a;
aud[30316]=16'h3a92;
aud[30317]=16'h3a89;
aud[30318]=16'h3a80;
aud[30319]=16'h3a78;
aud[30320]=16'h3a6f;
aud[30321]=16'h3a66;
aud[30322]=16'h3a5d;
aud[30323]=16'h3a54;
aud[30324]=16'h3a4c;
aud[30325]=16'h3a43;
aud[30326]=16'h3a3a;
aud[30327]=16'h3a31;
aud[30328]=16'h3a28;
aud[30329]=16'h3a1f;
aud[30330]=16'h3a16;
aud[30331]=16'h3a0d;
aud[30332]=16'h3a04;
aud[30333]=16'h39fb;
aud[30334]=16'h39f2;
aud[30335]=16'h39e9;
aud[30336]=16'h39e0;
aud[30337]=16'h39d6;
aud[30338]=16'h39cd;
aud[30339]=16'h39c4;
aud[30340]=16'h39bb;
aud[30341]=16'h39b1;
aud[30342]=16'h39a8;
aud[30343]=16'h399f;
aud[30344]=16'h3995;
aud[30345]=16'h398c;
aud[30346]=16'h3983;
aud[30347]=16'h3979;
aud[30348]=16'h3970;
aud[30349]=16'h3966;
aud[30350]=16'h395d;
aud[30351]=16'h3953;
aud[30352]=16'h394a;
aud[30353]=16'h3940;
aud[30354]=16'h3937;
aud[30355]=16'h392d;
aud[30356]=16'h3923;
aud[30357]=16'h391a;
aud[30358]=16'h3910;
aud[30359]=16'h3906;
aud[30360]=16'h38fd;
aud[30361]=16'h38f3;
aud[30362]=16'h38e9;
aud[30363]=16'h38df;
aud[30364]=16'h38d5;
aud[30365]=16'h38cb;
aud[30366]=16'h38c1;
aud[30367]=16'h38b8;
aud[30368]=16'h38ae;
aud[30369]=16'h38a4;
aud[30370]=16'h389a;
aud[30371]=16'h3890;
aud[30372]=16'h3886;
aud[30373]=16'h387b;
aud[30374]=16'h3871;
aud[30375]=16'h3867;
aud[30376]=16'h385d;
aud[30377]=16'h3853;
aud[30378]=16'h3849;
aud[30379]=16'h383f;
aud[30380]=16'h3834;
aud[30381]=16'h382a;
aud[30382]=16'h3820;
aud[30383]=16'h3815;
aud[30384]=16'h380b;
aud[30385]=16'h3801;
aud[30386]=16'h37f6;
aud[30387]=16'h37ec;
aud[30388]=16'h37e1;
aud[30389]=16'h37d7;
aud[30390]=16'h37cc;
aud[30391]=16'h37c2;
aud[30392]=16'h37b7;
aud[30393]=16'h37ad;
aud[30394]=16'h37a2;
aud[30395]=16'h3798;
aud[30396]=16'h378d;
aud[30397]=16'h3782;
aud[30398]=16'h3778;
aud[30399]=16'h376d;
aud[30400]=16'h3762;
aud[30401]=16'h3757;
aud[30402]=16'h374d;
aud[30403]=16'h3742;
aud[30404]=16'h3737;
aud[30405]=16'h372c;
aud[30406]=16'h3721;
aud[30407]=16'h3716;
aud[30408]=16'h370b;
aud[30409]=16'h3701;
aud[30410]=16'h36f6;
aud[30411]=16'h36eb;
aud[30412]=16'h36e0;
aud[30413]=16'h36d4;
aud[30414]=16'h36c9;
aud[30415]=16'h36be;
aud[30416]=16'h36b3;
aud[30417]=16'h36a8;
aud[30418]=16'h369d;
aud[30419]=16'h3692;
aud[30420]=16'h3686;
aud[30421]=16'h367b;
aud[30422]=16'h3670;
aud[30423]=16'h3665;
aud[30424]=16'h3659;
aud[30425]=16'h364e;
aud[30426]=16'h3643;
aud[30427]=16'h3637;
aud[30428]=16'h362c;
aud[30429]=16'h3620;
aud[30430]=16'h3615;
aud[30431]=16'h3609;
aud[30432]=16'h35fe;
aud[30433]=16'h35f2;
aud[30434]=16'h35e7;
aud[30435]=16'h35db;
aud[30436]=16'h35d0;
aud[30437]=16'h35c4;
aud[30438]=16'h35b8;
aud[30439]=16'h35ad;
aud[30440]=16'h35a1;
aud[30441]=16'h3595;
aud[30442]=16'h358a;
aud[30443]=16'h357e;
aud[30444]=16'h3572;
aud[30445]=16'h3566;
aud[30446]=16'h355a;
aud[30447]=16'h354f;
aud[30448]=16'h3543;
aud[30449]=16'h3537;
aud[30450]=16'h352b;
aud[30451]=16'h351f;
aud[30452]=16'h3513;
aud[30453]=16'h3507;
aud[30454]=16'h34fb;
aud[30455]=16'h34ef;
aud[30456]=16'h34e3;
aud[30457]=16'h34d7;
aud[30458]=16'h34cb;
aud[30459]=16'h34be;
aud[30460]=16'h34b2;
aud[30461]=16'h34a6;
aud[30462]=16'h349a;
aud[30463]=16'h348e;
aud[30464]=16'h3481;
aud[30465]=16'h3475;
aud[30466]=16'h3469;
aud[30467]=16'h345d;
aud[30468]=16'h3450;
aud[30469]=16'h3444;
aud[30470]=16'h3437;
aud[30471]=16'h342b;
aud[30472]=16'h341f;
aud[30473]=16'h3412;
aud[30474]=16'h3406;
aud[30475]=16'h33f9;
aud[30476]=16'h33ed;
aud[30477]=16'h33e0;
aud[30478]=16'h33d4;
aud[30479]=16'h33c7;
aud[30480]=16'h33ba;
aud[30481]=16'h33ae;
aud[30482]=16'h33a1;
aud[30483]=16'h3394;
aud[30484]=16'h3388;
aud[30485]=16'h337b;
aud[30486]=16'h336e;
aud[30487]=16'h3361;
aud[30488]=16'h3355;
aud[30489]=16'h3348;
aud[30490]=16'h333b;
aud[30491]=16'h332e;
aud[30492]=16'h3321;
aud[30493]=16'h3314;
aud[30494]=16'h3307;
aud[30495]=16'h32fa;
aud[30496]=16'h32ed;
aud[30497]=16'h32e0;
aud[30498]=16'h32d3;
aud[30499]=16'h32c6;
aud[30500]=16'h32b9;
aud[30501]=16'h32ac;
aud[30502]=16'h329f;
aud[30503]=16'h3292;
aud[30504]=16'h3285;
aud[30505]=16'h3278;
aud[30506]=16'h326a;
aud[30507]=16'h325d;
aud[30508]=16'h3250;
aud[30509]=16'h3243;
aud[30510]=16'h3235;
aud[30511]=16'h3228;
aud[30512]=16'h321b;
aud[30513]=16'h320d;
aud[30514]=16'h3200;
aud[30515]=16'h31f3;
aud[30516]=16'h31e5;
aud[30517]=16'h31d8;
aud[30518]=16'h31ca;
aud[30519]=16'h31bd;
aud[30520]=16'h31af;
aud[30521]=16'h31a2;
aud[30522]=16'h3194;
aud[30523]=16'h3187;
aud[30524]=16'h3179;
aud[30525]=16'h316b;
aud[30526]=16'h315e;
aud[30527]=16'h3150;
aud[30528]=16'h3142;
aud[30529]=16'h3135;
aud[30530]=16'h3127;
aud[30531]=16'h3119;
aud[30532]=16'h310b;
aud[30533]=16'h30fe;
aud[30534]=16'h30f0;
aud[30535]=16'h30e2;
aud[30536]=16'h30d4;
aud[30537]=16'h30c6;
aud[30538]=16'h30b8;
aud[30539]=16'h30aa;
aud[30540]=16'h309d;
aud[30541]=16'h308f;
aud[30542]=16'h3081;
aud[30543]=16'h3073;
aud[30544]=16'h3065;
aud[30545]=16'h3057;
aud[30546]=16'h3048;
aud[30547]=16'h303a;
aud[30548]=16'h302c;
aud[30549]=16'h301e;
aud[30550]=16'h3010;
aud[30551]=16'h3002;
aud[30552]=16'h2ff4;
aud[30553]=16'h2fe5;
aud[30554]=16'h2fd7;
aud[30555]=16'h2fc9;
aud[30556]=16'h2fbb;
aud[30557]=16'h2fac;
aud[30558]=16'h2f9e;
aud[30559]=16'h2f90;
aud[30560]=16'h2f81;
aud[30561]=16'h2f73;
aud[30562]=16'h2f65;
aud[30563]=16'h2f56;
aud[30564]=16'h2f48;
aud[30565]=16'h2f39;
aud[30566]=16'h2f2b;
aud[30567]=16'h2f1c;
aud[30568]=16'h2f0e;
aud[30569]=16'h2eff;
aud[30570]=16'h2ef1;
aud[30571]=16'h2ee2;
aud[30572]=16'h2ed3;
aud[30573]=16'h2ec5;
aud[30574]=16'h2eb6;
aud[30575]=16'h2ea7;
aud[30576]=16'h2e99;
aud[30577]=16'h2e8a;
aud[30578]=16'h2e7b;
aud[30579]=16'h2e6d;
aud[30580]=16'h2e5e;
aud[30581]=16'h2e4f;
aud[30582]=16'h2e40;
aud[30583]=16'h2e31;
aud[30584]=16'h2e22;
aud[30585]=16'h2e14;
aud[30586]=16'h2e05;
aud[30587]=16'h2df6;
aud[30588]=16'h2de7;
aud[30589]=16'h2dd8;
aud[30590]=16'h2dc9;
aud[30591]=16'h2dba;
aud[30592]=16'h2dab;
aud[30593]=16'h2d9c;
aud[30594]=16'h2d8d;
aud[30595]=16'h2d7e;
aud[30596]=16'h2d6f;
aud[30597]=16'h2d60;
aud[30598]=16'h2d50;
aud[30599]=16'h2d41;
aud[30600]=16'h2d32;
aud[30601]=16'h2d23;
aud[30602]=16'h2d14;
aud[30603]=16'h2d04;
aud[30604]=16'h2cf5;
aud[30605]=16'h2ce6;
aud[30606]=16'h2cd7;
aud[30607]=16'h2cc7;
aud[30608]=16'h2cb8;
aud[30609]=16'h2ca9;
aud[30610]=16'h2c99;
aud[30611]=16'h2c8a;
aud[30612]=16'h2c7a;
aud[30613]=16'h2c6b;
aud[30614]=16'h2c5c;
aud[30615]=16'h2c4c;
aud[30616]=16'h2c3d;
aud[30617]=16'h2c2d;
aud[30618]=16'h2c1e;
aud[30619]=16'h2c0e;
aud[30620]=16'h2bfe;
aud[30621]=16'h2bef;
aud[30622]=16'h2bdf;
aud[30623]=16'h2bd0;
aud[30624]=16'h2bc0;
aud[30625]=16'h2bb0;
aud[30626]=16'h2ba1;
aud[30627]=16'h2b91;
aud[30628]=16'h2b81;
aud[30629]=16'h2b71;
aud[30630]=16'h2b62;
aud[30631]=16'h2b52;
aud[30632]=16'h2b42;
aud[30633]=16'h2b32;
aud[30634]=16'h2b22;
aud[30635]=16'h2b13;
aud[30636]=16'h2b03;
aud[30637]=16'h2af3;
aud[30638]=16'h2ae3;
aud[30639]=16'h2ad3;
aud[30640]=16'h2ac3;
aud[30641]=16'h2ab3;
aud[30642]=16'h2aa3;
aud[30643]=16'h2a93;
aud[30644]=16'h2a83;
aud[30645]=16'h2a73;
aud[30646]=16'h2a63;
aud[30647]=16'h2a53;
aud[30648]=16'h2a43;
aud[30649]=16'h2a33;
aud[30650]=16'h2a23;
aud[30651]=16'h2a12;
aud[30652]=16'h2a02;
aud[30653]=16'h29f2;
aud[30654]=16'h29e2;
aud[30655]=16'h29d2;
aud[30656]=16'h29c1;
aud[30657]=16'h29b1;
aud[30658]=16'h29a1;
aud[30659]=16'h2991;
aud[30660]=16'h2980;
aud[30661]=16'h2970;
aud[30662]=16'h2960;
aud[30663]=16'h294f;
aud[30664]=16'h293f;
aud[30665]=16'h292e;
aud[30666]=16'h291e;
aud[30667]=16'h290e;
aud[30668]=16'h28fd;
aud[30669]=16'h28ed;
aud[30670]=16'h28dc;
aud[30671]=16'h28cc;
aud[30672]=16'h28bb;
aud[30673]=16'h28aa;
aud[30674]=16'h289a;
aud[30675]=16'h2889;
aud[30676]=16'h2879;
aud[30677]=16'h2868;
aud[30678]=16'h2857;
aud[30679]=16'h2847;
aud[30680]=16'h2836;
aud[30681]=16'h2825;
aud[30682]=16'h2815;
aud[30683]=16'h2804;
aud[30684]=16'h27f3;
aud[30685]=16'h27e2;
aud[30686]=16'h27d2;
aud[30687]=16'h27c1;
aud[30688]=16'h27b0;
aud[30689]=16'h279f;
aud[30690]=16'h278e;
aud[30691]=16'h277e;
aud[30692]=16'h276d;
aud[30693]=16'h275c;
aud[30694]=16'h274b;
aud[30695]=16'h273a;
aud[30696]=16'h2729;
aud[30697]=16'h2718;
aud[30698]=16'h2707;
aud[30699]=16'h26f6;
aud[30700]=16'h26e5;
aud[30701]=16'h26d4;
aud[30702]=16'h26c3;
aud[30703]=16'h26b2;
aud[30704]=16'h26a1;
aud[30705]=16'h2690;
aud[30706]=16'h267e;
aud[30707]=16'h266d;
aud[30708]=16'h265c;
aud[30709]=16'h264b;
aud[30710]=16'h263a;
aud[30711]=16'h2629;
aud[30712]=16'h2617;
aud[30713]=16'h2606;
aud[30714]=16'h25f5;
aud[30715]=16'h25e4;
aud[30716]=16'h25d2;
aud[30717]=16'h25c1;
aud[30718]=16'h25b0;
aud[30719]=16'h259e;
aud[30720]=16'h258d;
aud[30721]=16'h257c;
aud[30722]=16'h256a;
aud[30723]=16'h2559;
aud[30724]=16'h2547;
aud[30725]=16'h2536;
aud[30726]=16'h2524;
aud[30727]=16'h2513;
aud[30728]=16'h2501;
aud[30729]=16'h24f0;
aud[30730]=16'h24de;
aud[30731]=16'h24cd;
aud[30732]=16'h24bb;
aud[30733]=16'h24aa;
aud[30734]=16'h2498;
aud[30735]=16'h2487;
aud[30736]=16'h2475;
aud[30737]=16'h2463;
aud[30738]=16'h2452;
aud[30739]=16'h2440;
aud[30740]=16'h242e;
aud[30741]=16'h241d;
aud[30742]=16'h240b;
aud[30743]=16'h23f9;
aud[30744]=16'h23e7;
aud[30745]=16'h23d6;
aud[30746]=16'h23c4;
aud[30747]=16'h23b2;
aud[30748]=16'h23a0;
aud[30749]=16'h238e;
aud[30750]=16'h237d;
aud[30751]=16'h236b;
aud[30752]=16'h2359;
aud[30753]=16'h2347;
aud[30754]=16'h2335;
aud[30755]=16'h2323;
aud[30756]=16'h2311;
aud[30757]=16'h22ff;
aud[30758]=16'h22ed;
aud[30759]=16'h22db;
aud[30760]=16'h22c9;
aud[30761]=16'h22b7;
aud[30762]=16'h22a5;
aud[30763]=16'h2293;
aud[30764]=16'h2281;
aud[30765]=16'h226f;
aud[30766]=16'h225d;
aud[30767]=16'h224b;
aud[30768]=16'h2239;
aud[30769]=16'h2227;
aud[30770]=16'h2215;
aud[30771]=16'h2202;
aud[30772]=16'h21f0;
aud[30773]=16'h21de;
aud[30774]=16'h21cc;
aud[30775]=16'h21ba;
aud[30776]=16'h21a7;
aud[30777]=16'h2195;
aud[30778]=16'h2183;
aud[30779]=16'h2171;
aud[30780]=16'h215e;
aud[30781]=16'h214c;
aud[30782]=16'h213a;
aud[30783]=16'h2127;
aud[30784]=16'h2115;
aud[30785]=16'h2103;
aud[30786]=16'h20f0;
aud[30787]=16'h20de;
aud[30788]=16'h20cb;
aud[30789]=16'h20b9;
aud[30790]=16'h20a7;
aud[30791]=16'h2094;
aud[30792]=16'h2082;
aud[30793]=16'h206f;
aud[30794]=16'h205d;
aud[30795]=16'h204a;
aud[30796]=16'h2038;
aud[30797]=16'h2025;
aud[30798]=16'h2013;
aud[30799]=16'h2000;
aud[30800]=16'h1fed;
aud[30801]=16'h1fdb;
aud[30802]=16'h1fc8;
aud[30803]=16'h1fb6;
aud[30804]=16'h1fa3;
aud[30805]=16'h1f90;
aud[30806]=16'h1f7e;
aud[30807]=16'h1f6b;
aud[30808]=16'h1f58;
aud[30809]=16'h1f46;
aud[30810]=16'h1f33;
aud[30811]=16'h1f20;
aud[30812]=16'h1f0d;
aud[30813]=16'h1efb;
aud[30814]=16'h1ee8;
aud[30815]=16'h1ed5;
aud[30816]=16'h1ec2;
aud[30817]=16'h1eaf;
aud[30818]=16'h1e9d;
aud[30819]=16'h1e8a;
aud[30820]=16'h1e77;
aud[30821]=16'h1e64;
aud[30822]=16'h1e51;
aud[30823]=16'h1e3e;
aud[30824]=16'h1e2b;
aud[30825]=16'h1e18;
aud[30826]=16'h1e06;
aud[30827]=16'h1df3;
aud[30828]=16'h1de0;
aud[30829]=16'h1dcd;
aud[30830]=16'h1dba;
aud[30831]=16'h1da7;
aud[30832]=16'h1d94;
aud[30833]=16'h1d81;
aud[30834]=16'h1d6e;
aud[30835]=16'h1d5b;
aud[30836]=16'h1d47;
aud[30837]=16'h1d34;
aud[30838]=16'h1d21;
aud[30839]=16'h1d0e;
aud[30840]=16'h1cfb;
aud[30841]=16'h1ce8;
aud[30842]=16'h1cd5;
aud[30843]=16'h1cc2;
aud[30844]=16'h1cae;
aud[30845]=16'h1c9b;
aud[30846]=16'h1c88;
aud[30847]=16'h1c75;
aud[30848]=16'h1c62;
aud[30849]=16'h1c4e;
aud[30850]=16'h1c3b;
aud[30851]=16'h1c28;
aud[30852]=16'h1c15;
aud[30853]=16'h1c01;
aud[30854]=16'h1bee;
aud[30855]=16'h1bdb;
aud[30856]=16'h1bc8;
aud[30857]=16'h1bb4;
aud[30858]=16'h1ba1;
aud[30859]=16'h1b8d;
aud[30860]=16'h1b7a;
aud[30861]=16'h1b67;
aud[30862]=16'h1b53;
aud[30863]=16'h1b40;
aud[30864]=16'h1b2d;
aud[30865]=16'h1b19;
aud[30866]=16'h1b06;
aud[30867]=16'h1af2;
aud[30868]=16'h1adf;
aud[30869]=16'h1acb;
aud[30870]=16'h1ab8;
aud[30871]=16'h1aa4;
aud[30872]=16'h1a91;
aud[30873]=16'h1a7d;
aud[30874]=16'h1a6a;
aud[30875]=16'h1a56;
aud[30876]=16'h1a43;
aud[30877]=16'h1a2f;
aud[30878]=16'h1a1c;
aud[30879]=16'h1a08;
aud[30880]=16'h19f4;
aud[30881]=16'h19e1;
aud[30882]=16'h19cd;
aud[30883]=16'h19ba;
aud[30884]=16'h19a6;
aud[30885]=16'h1992;
aud[30886]=16'h197f;
aud[30887]=16'h196b;
aud[30888]=16'h1957;
aud[30889]=16'h1943;
aud[30890]=16'h1930;
aud[30891]=16'h191c;
aud[30892]=16'h1908;
aud[30893]=16'h18f5;
aud[30894]=16'h18e1;
aud[30895]=16'h18cd;
aud[30896]=16'h18b9;
aud[30897]=16'h18a5;
aud[30898]=16'h1892;
aud[30899]=16'h187e;
aud[30900]=16'h186a;
aud[30901]=16'h1856;
aud[30902]=16'h1842;
aud[30903]=16'h182f;
aud[30904]=16'h181b;
aud[30905]=16'h1807;
aud[30906]=16'h17f3;
aud[30907]=16'h17df;
aud[30908]=16'h17cb;
aud[30909]=16'h17b7;
aud[30910]=16'h17a3;
aud[30911]=16'h178f;
aud[30912]=16'h177b;
aud[30913]=16'h1767;
aud[30914]=16'h1753;
aud[30915]=16'h1740;
aud[30916]=16'h172c;
aud[30917]=16'h1718;
aud[30918]=16'h1704;
aud[30919]=16'h16f0;
aud[30920]=16'h16db;
aud[30921]=16'h16c7;
aud[30922]=16'h16b3;
aud[30923]=16'h169f;
aud[30924]=16'h168b;
aud[30925]=16'h1677;
aud[30926]=16'h1663;
aud[30927]=16'h164f;
aud[30928]=16'h163b;
aud[30929]=16'h1627;
aud[30930]=16'h1613;
aud[30931]=16'h15ff;
aud[30932]=16'h15ea;
aud[30933]=16'h15d6;
aud[30934]=16'h15c2;
aud[30935]=16'h15ae;
aud[30936]=16'h159a;
aud[30937]=16'h1586;
aud[30938]=16'h1571;
aud[30939]=16'h155d;
aud[30940]=16'h1549;
aud[30941]=16'h1535;
aud[30942]=16'h1520;
aud[30943]=16'h150c;
aud[30944]=16'h14f8;
aud[30945]=16'h14e4;
aud[30946]=16'h14cf;
aud[30947]=16'h14bb;
aud[30948]=16'h14a7;
aud[30949]=16'h1492;
aud[30950]=16'h147e;
aud[30951]=16'h146a;
aud[30952]=16'h1455;
aud[30953]=16'h1441;
aud[30954]=16'h142d;
aud[30955]=16'h1418;
aud[30956]=16'h1404;
aud[30957]=16'h13f0;
aud[30958]=16'h13db;
aud[30959]=16'h13c7;
aud[30960]=16'h13b3;
aud[30961]=16'h139e;
aud[30962]=16'h138a;
aud[30963]=16'h1375;
aud[30964]=16'h1361;
aud[30965]=16'h134c;
aud[30966]=16'h1338;
aud[30967]=16'h1323;
aud[30968]=16'h130f;
aud[30969]=16'h12fb;
aud[30970]=16'h12e6;
aud[30971]=16'h12d2;
aud[30972]=16'h12bd;
aud[30973]=16'h12a9;
aud[30974]=16'h1294;
aud[30975]=16'h127f;
aud[30976]=16'h126b;
aud[30977]=16'h1256;
aud[30978]=16'h1242;
aud[30979]=16'h122d;
aud[30980]=16'h1219;
aud[30981]=16'h1204;
aud[30982]=16'h11f0;
aud[30983]=16'h11db;
aud[30984]=16'h11c6;
aud[30985]=16'h11b2;
aud[30986]=16'h119d;
aud[30987]=16'h1189;
aud[30988]=16'h1174;
aud[30989]=16'h115f;
aud[30990]=16'h114b;
aud[30991]=16'h1136;
aud[30992]=16'h1121;
aud[30993]=16'h110d;
aud[30994]=16'h10f8;
aud[30995]=16'h10e3;
aud[30996]=16'h10cf;
aud[30997]=16'h10ba;
aud[30998]=16'h10a5;
aud[30999]=16'h1090;
aud[31000]=16'h107c;
aud[31001]=16'h1067;
aud[31002]=16'h1052;
aud[31003]=16'h103e;
aud[31004]=16'h1029;
aud[31005]=16'h1014;
aud[31006]=16'hfff;
aud[31007]=16'hfeb;
aud[31008]=16'hfd6;
aud[31009]=16'hfc1;
aud[31010]=16'hfac;
aud[31011]=16'hf97;
aud[31012]=16'hf83;
aud[31013]=16'hf6e;
aud[31014]=16'hf59;
aud[31015]=16'hf44;
aud[31016]=16'hf2f;
aud[31017]=16'hf1a;
aud[31018]=16'hf06;
aud[31019]=16'hef1;
aud[31020]=16'hedc;
aud[31021]=16'hec7;
aud[31022]=16'heb2;
aud[31023]=16'he9d;
aud[31024]=16'he88;
aud[31025]=16'he74;
aud[31026]=16'he5f;
aud[31027]=16'he4a;
aud[31028]=16'he35;
aud[31029]=16'he20;
aud[31030]=16'he0b;
aud[31031]=16'hdf6;
aud[31032]=16'hde1;
aud[31033]=16'hdcc;
aud[31034]=16'hdb7;
aud[31035]=16'hda2;
aud[31036]=16'hd8d;
aud[31037]=16'hd78;
aud[31038]=16'hd63;
aud[31039]=16'hd4e;
aud[31040]=16'hd39;
aud[31041]=16'hd24;
aud[31042]=16'hd0f;
aud[31043]=16'hcfa;
aud[31044]=16'hce5;
aud[31045]=16'hcd0;
aud[31046]=16'hcbb;
aud[31047]=16'hca6;
aud[31048]=16'hc91;
aud[31049]=16'hc7c;
aud[31050]=16'hc67;
aud[31051]=16'hc52;
aud[31052]=16'hc3d;
aud[31053]=16'hc28;
aud[31054]=16'hc13;
aud[31055]=16'hbfe;
aud[31056]=16'hbe9;
aud[31057]=16'hbd4;
aud[31058]=16'hbbf;
aud[31059]=16'hbaa;
aud[31060]=16'hb95;
aud[31061]=16'hb80;
aud[31062]=16'hb6a;
aud[31063]=16'hb55;
aud[31064]=16'hb40;
aud[31065]=16'hb2b;
aud[31066]=16'hb16;
aud[31067]=16'hb01;
aud[31068]=16'haec;
aud[31069]=16'had7;
aud[31070]=16'hac1;
aud[31071]=16'haac;
aud[31072]=16'ha97;
aud[31073]=16'ha82;
aud[31074]=16'ha6d;
aud[31075]=16'ha58;
aud[31076]=16'ha43;
aud[31077]=16'ha2d;
aud[31078]=16'ha18;
aud[31079]=16'ha03;
aud[31080]=16'h9ee;
aud[31081]=16'h9d9;
aud[31082]=16'h9c3;
aud[31083]=16'h9ae;
aud[31084]=16'h999;
aud[31085]=16'h984;
aud[31086]=16'h96f;
aud[31087]=16'h959;
aud[31088]=16'h944;
aud[31089]=16'h92f;
aud[31090]=16'h91a;
aud[31091]=16'h905;
aud[31092]=16'h8ef;
aud[31093]=16'h8da;
aud[31094]=16'h8c5;
aud[31095]=16'h8b0;
aud[31096]=16'h89a;
aud[31097]=16'h885;
aud[31098]=16'h870;
aud[31099]=16'h85b;
aud[31100]=16'h845;
aud[31101]=16'h830;
aud[31102]=16'h81b;
aud[31103]=16'h805;
aud[31104]=16'h7f0;
aud[31105]=16'h7db;
aud[31106]=16'h7c6;
aud[31107]=16'h7b0;
aud[31108]=16'h79b;
aud[31109]=16'h786;
aud[31110]=16'h770;
aud[31111]=16'h75b;
aud[31112]=16'h746;
aud[31113]=16'h731;
aud[31114]=16'h71b;
aud[31115]=16'h706;
aud[31116]=16'h6f1;
aud[31117]=16'h6db;
aud[31118]=16'h6c6;
aud[31119]=16'h6b1;
aud[31120]=16'h69b;
aud[31121]=16'h686;
aud[31122]=16'h671;
aud[31123]=16'h65b;
aud[31124]=16'h646;
aud[31125]=16'h631;
aud[31126]=16'h61b;
aud[31127]=16'h606;
aud[31128]=16'h5f1;
aud[31129]=16'h5db;
aud[31130]=16'h5c6;
aud[31131]=16'h5b0;
aud[31132]=16'h59b;
aud[31133]=16'h586;
aud[31134]=16'h570;
aud[31135]=16'h55b;
aud[31136]=16'h546;
aud[31137]=16'h530;
aud[31138]=16'h51b;
aud[31139]=16'h505;
aud[31140]=16'h4f0;
aud[31141]=16'h4db;
aud[31142]=16'h4c5;
aud[31143]=16'h4b0;
aud[31144]=16'h49b;
aud[31145]=16'h485;
aud[31146]=16'h470;
aud[31147]=16'h45a;
aud[31148]=16'h445;
aud[31149]=16'h430;
aud[31150]=16'h41a;
aud[31151]=16'h405;
aud[31152]=16'h3ef;
aud[31153]=16'h3da;
aud[31154]=16'h3c5;
aud[31155]=16'h3af;
aud[31156]=16'h39a;
aud[31157]=16'h384;
aud[31158]=16'h36f;
aud[31159]=16'h359;
aud[31160]=16'h344;
aud[31161]=16'h32f;
aud[31162]=16'h319;
aud[31163]=16'h304;
aud[31164]=16'h2ee;
aud[31165]=16'h2d9;
aud[31166]=16'h2c4;
aud[31167]=16'h2ae;
aud[31168]=16'h299;
aud[31169]=16'h283;
aud[31170]=16'h26e;
aud[31171]=16'h258;
aud[31172]=16'h243;
aud[31173]=16'h22e;
aud[31174]=16'h218;
aud[31175]=16'h203;
aud[31176]=16'h1ed;
aud[31177]=16'h1d8;
aud[31178]=16'h1c2;
aud[31179]=16'h1ad;
aud[31180]=16'h197;
aud[31181]=16'h182;
aud[31182]=16'h16d;
aud[31183]=16'h157;
aud[31184]=16'h142;
aud[31185]=16'h12c;
aud[31186]=16'h117;
aud[31187]=16'h101;
aud[31188]=16'hec;
aud[31189]=16'hd6;
aud[31190]=16'hc1;
aud[31191]=16'hac;
aud[31192]=16'h96;
aud[31193]=16'h81;
aud[31194]=16'h6b;
aud[31195]=16'h56;
aud[31196]=16'h40;
aud[31197]=16'h2b;
aud[31198]=16'h15;
aud[31199]=16'h0;
aud[31200]=16'hffeb;
aud[31201]=16'hffd5;
aud[31202]=16'hffc0;
aud[31203]=16'hffaa;
aud[31204]=16'hff95;
aud[31205]=16'hff7f;
aud[31206]=16'hff6a;
aud[31207]=16'hff54;
aud[31208]=16'hff3f;
aud[31209]=16'hff2a;
aud[31210]=16'hff14;
aud[31211]=16'hfeff;
aud[31212]=16'hfee9;
aud[31213]=16'hfed4;
aud[31214]=16'hfebe;
aud[31215]=16'hfea9;
aud[31216]=16'hfe93;
aud[31217]=16'hfe7e;
aud[31218]=16'hfe69;
aud[31219]=16'hfe53;
aud[31220]=16'hfe3e;
aud[31221]=16'hfe28;
aud[31222]=16'hfe13;
aud[31223]=16'hfdfd;
aud[31224]=16'hfde8;
aud[31225]=16'hfdd2;
aud[31226]=16'hfdbd;
aud[31227]=16'hfda8;
aud[31228]=16'hfd92;
aud[31229]=16'hfd7d;
aud[31230]=16'hfd67;
aud[31231]=16'hfd52;
aud[31232]=16'hfd3c;
aud[31233]=16'hfd27;
aud[31234]=16'hfd12;
aud[31235]=16'hfcfc;
aud[31236]=16'hfce7;
aud[31237]=16'hfcd1;
aud[31238]=16'hfcbc;
aud[31239]=16'hfca7;
aud[31240]=16'hfc91;
aud[31241]=16'hfc7c;
aud[31242]=16'hfc66;
aud[31243]=16'hfc51;
aud[31244]=16'hfc3b;
aud[31245]=16'hfc26;
aud[31246]=16'hfc11;
aud[31247]=16'hfbfb;
aud[31248]=16'hfbe6;
aud[31249]=16'hfbd0;
aud[31250]=16'hfbbb;
aud[31251]=16'hfba6;
aud[31252]=16'hfb90;
aud[31253]=16'hfb7b;
aud[31254]=16'hfb65;
aud[31255]=16'hfb50;
aud[31256]=16'hfb3b;
aud[31257]=16'hfb25;
aud[31258]=16'hfb10;
aud[31259]=16'hfafb;
aud[31260]=16'hfae5;
aud[31261]=16'hfad0;
aud[31262]=16'hfaba;
aud[31263]=16'hfaa5;
aud[31264]=16'hfa90;
aud[31265]=16'hfa7a;
aud[31266]=16'hfa65;
aud[31267]=16'hfa50;
aud[31268]=16'hfa3a;
aud[31269]=16'hfa25;
aud[31270]=16'hfa0f;
aud[31271]=16'hf9fa;
aud[31272]=16'hf9e5;
aud[31273]=16'hf9cf;
aud[31274]=16'hf9ba;
aud[31275]=16'hf9a5;
aud[31276]=16'hf98f;
aud[31277]=16'hf97a;
aud[31278]=16'hf965;
aud[31279]=16'hf94f;
aud[31280]=16'hf93a;
aud[31281]=16'hf925;
aud[31282]=16'hf90f;
aud[31283]=16'hf8fa;
aud[31284]=16'hf8e5;
aud[31285]=16'hf8cf;
aud[31286]=16'hf8ba;
aud[31287]=16'hf8a5;
aud[31288]=16'hf890;
aud[31289]=16'hf87a;
aud[31290]=16'hf865;
aud[31291]=16'hf850;
aud[31292]=16'hf83a;
aud[31293]=16'hf825;
aud[31294]=16'hf810;
aud[31295]=16'hf7fb;
aud[31296]=16'hf7e5;
aud[31297]=16'hf7d0;
aud[31298]=16'hf7bb;
aud[31299]=16'hf7a5;
aud[31300]=16'hf790;
aud[31301]=16'hf77b;
aud[31302]=16'hf766;
aud[31303]=16'hf750;
aud[31304]=16'hf73b;
aud[31305]=16'hf726;
aud[31306]=16'hf711;
aud[31307]=16'hf6fb;
aud[31308]=16'hf6e6;
aud[31309]=16'hf6d1;
aud[31310]=16'hf6bc;
aud[31311]=16'hf6a7;
aud[31312]=16'hf691;
aud[31313]=16'hf67c;
aud[31314]=16'hf667;
aud[31315]=16'hf652;
aud[31316]=16'hf63d;
aud[31317]=16'hf627;
aud[31318]=16'hf612;
aud[31319]=16'hf5fd;
aud[31320]=16'hf5e8;
aud[31321]=16'hf5d3;
aud[31322]=16'hf5bd;
aud[31323]=16'hf5a8;
aud[31324]=16'hf593;
aud[31325]=16'hf57e;
aud[31326]=16'hf569;
aud[31327]=16'hf554;
aud[31328]=16'hf53f;
aud[31329]=16'hf529;
aud[31330]=16'hf514;
aud[31331]=16'hf4ff;
aud[31332]=16'hf4ea;
aud[31333]=16'hf4d5;
aud[31334]=16'hf4c0;
aud[31335]=16'hf4ab;
aud[31336]=16'hf496;
aud[31337]=16'hf480;
aud[31338]=16'hf46b;
aud[31339]=16'hf456;
aud[31340]=16'hf441;
aud[31341]=16'hf42c;
aud[31342]=16'hf417;
aud[31343]=16'hf402;
aud[31344]=16'hf3ed;
aud[31345]=16'hf3d8;
aud[31346]=16'hf3c3;
aud[31347]=16'hf3ae;
aud[31348]=16'hf399;
aud[31349]=16'hf384;
aud[31350]=16'hf36f;
aud[31351]=16'hf35a;
aud[31352]=16'hf345;
aud[31353]=16'hf330;
aud[31354]=16'hf31b;
aud[31355]=16'hf306;
aud[31356]=16'hf2f1;
aud[31357]=16'hf2dc;
aud[31358]=16'hf2c7;
aud[31359]=16'hf2b2;
aud[31360]=16'hf29d;
aud[31361]=16'hf288;
aud[31362]=16'hf273;
aud[31363]=16'hf25e;
aud[31364]=16'hf249;
aud[31365]=16'hf234;
aud[31366]=16'hf21f;
aud[31367]=16'hf20a;
aud[31368]=16'hf1f5;
aud[31369]=16'hf1e0;
aud[31370]=16'hf1cb;
aud[31371]=16'hf1b6;
aud[31372]=16'hf1a1;
aud[31373]=16'hf18c;
aud[31374]=16'hf178;
aud[31375]=16'hf163;
aud[31376]=16'hf14e;
aud[31377]=16'hf139;
aud[31378]=16'hf124;
aud[31379]=16'hf10f;
aud[31380]=16'hf0fa;
aud[31381]=16'hf0e6;
aud[31382]=16'hf0d1;
aud[31383]=16'hf0bc;
aud[31384]=16'hf0a7;
aud[31385]=16'hf092;
aud[31386]=16'hf07d;
aud[31387]=16'hf069;
aud[31388]=16'hf054;
aud[31389]=16'hf03f;
aud[31390]=16'hf02a;
aud[31391]=16'hf015;
aud[31392]=16'hf001;
aud[31393]=16'hefec;
aud[31394]=16'hefd7;
aud[31395]=16'hefc2;
aud[31396]=16'hefae;
aud[31397]=16'hef99;
aud[31398]=16'hef84;
aud[31399]=16'hef70;
aud[31400]=16'hef5b;
aud[31401]=16'hef46;
aud[31402]=16'hef31;
aud[31403]=16'hef1d;
aud[31404]=16'hef08;
aud[31405]=16'heef3;
aud[31406]=16'heedf;
aud[31407]=16'heeca;
aud[31408]=16'heeb5;
aud[31409]=16'heea1;
aud[31410]=16'hee8c;
aud[31411]=16'hee77;
aud[31412]=16'hee63;
aud[31413]=16'hee4e;
aud[31414]=16'hee3a;
aud[31415]=16'hee25;
aud[31416]=16'hee10;
aud[31417]=16'hedfc;
aud[31418]=16'hede7;
aud[31419]=16'hedd3;
aud[31420]=16'hedbe;
aud[31421]=16'hedaa;
aud[31422]=16'hed95;
aud[31423]=16'hed81;
aud[31424]=16'hed6c;
aud[31425]=16'hed57;
aud[31426]=16'hed43;
aud[31427]=16'hed2e;
aud[31428]=16'hed1a;
aud[31429]=16'hed05;
aud[31430]=16'hecf1;
aud[31431]=16'hecdd;
aud[31432]=16'hecc8;
aud[31433]=16'hecb4;
aud[31434]=16'hec9f;
aud[31435]=16'hec8b;
aud[31436]=16'hec76;
aud[31437]=16'hec62;
aud[31438]=16'hec4d;
aud[31439]=16'hec39;
aud[31440]=16'hec25;
aud[31441]=16'hec10;
aud[31442]=16'hebfc;
aud[31443]=16'hebe8;
aud[31444]=16'hebd3;
aud[31445]=16'hebbf;
aud[31446]=16'hebab;
aud[31447]=16'heb96;
aud[31448]=16'heb82;
aud[31449]=16'heb6e;
aud[31450]=16'heb59;
aud[31451]=16'heb45;
aud[31452]=16'heb31;
aud[31453]=16'heb1c;
aud[31454]=16'heb08;
aud[31455]=16'heaf4;
aud[31456]=16'heae0;
aud[31457]=16'heacb;
aud[31458]=16'heab7;
aud[31459]=16'heaa3;
aud[31460]=16'hea8f;
aud[31461]=16'hea7a;
aud[31462]=16'hea66;
aud[31463]=16'hea52;
aud[31464]=16'hea3e;
aud[31465]=16'hea2a;
aud[31466]=16'hea16;
aud[31467]=16'hea01;
aud[31468]=16'he9ed;
aud[31469]=16'he9d9;
aud[31470]=16'he9c5;
aud[31471]=16'he9b1;
aud[31472]=16'he99d;
aud[31473]=16'he989;
aud[31474]=16'he975;
aud[31475]=16'he961;
aud[31476]=16'he94d;
aud[31477]=16'he939;
aud[31478]=16'he925;
aud[31479]=16'he910;
aud[31480]=16'he8fc;
aud[31481]=16'he8e8;
aud[31482]=16'he8d4;
aud[31483]=16'he8c0;
aud[31484]=16'he8ad;
aud[31485]=16'he899;
aud[31486]=16'he885;
aud[31487]=16'he871;
aud[31488]=16'he85d;
aud[31489]=16'he849;
aud[31490]=16'he835;
aud[31491]=16'he821;
aud[31492]=16'he80d;
aud[31493]=16'he7f9;
aud[31494]=16'he7e5;
aud[31495]=16'he7d1;
aud[31496]=16'he7be;
aud[31497]=16'he7aa;
aud[31498]=16'he796;
aud[31499]=16'he782;
aud[31500]=16'he76e;
aud[31501]=16'he75b;
aud[31502]=16'he747;
aud[31503]=16'he733;
aud[31504]=16'he71f;
aud[31505]=16'he70b;
aud[31506]=16'he6f8;
aud[31507]=16'he6e4;
aud[31508]=16'he6d0;
aud[31509]=16'he6bd;
aud[31510]=16'he6a9;
aud[31511]=16'he695;
aud[31512]=16'he681;
aud[31513]=16'he66e;
aud[31514]=16'he65a;
aud[31515]=16'he646;
aud[31516]=16'he633;
aud[31517]=16'he61f;
aud[31518]=16'he60c;
aud[31519]=16'he5f8;
aud[31520]=16'he5e4;
aud[31521]=16'he5d1;
aud[31522]=16'he5bd;
aud[31523]=16'he5aa;
aud[31524]=16'he596;
aud[31525]=16'he583;
aud[31526]=16'he56f;
aud[31527]=16'he55c;
aud[31528]=16'he548;
aud[31529]=16'he535;
aud[31530]=16'he521;
aud[31531]=16'he50e;
aud[31532]=16'he4fa;
aud[31533]=16'he4e7;
aud[31534]=16'he4d3;
aud[31535]=16'he4c0;
aud[31536]=16'he4ad;
aud[31537]=16'he499;
aud[31538]=16'he486;
aud[31539]=16'he473;
aud[31540]=16'he45f;
aud[31541]=16'he44c;
aud[31542]=16'he438;
aud[31543]=16'he425;
aud[31544]=16'he412;
aud[31545]=16'he3ff;
aud[31546]=16'he3eb;
aud[31547]=16'he3d8;
aud[31548]=16'he3c5;
aud[31549]=16'he3b2;
aud[31550]=16'he39e;
aud[31551]=16'he38b;
aud[31552]=16'he378;
aud[31553]=16'he365;
aud[31554]=16'he352;
aud[31555]=16'he33e;
aud[31556]=16'he32b;
aud[31557]=16'he318;
aud[31558]=16'he305;
aud[31559]=16'he2f2;
aud[31560]=16'he2df;
aud[31561]=16'he2cc;
aud[31562]=16'he2b9;
aud[31563]=16'he2a5;
aud[31564]=16'he292;
aud[31565]=16'he27f;
aud[31566]=16'he26c;
aud[31567]=16'he259;
aud[31568]=16'he246;
aud[31569]=16'he233;
aud[31570]=16'he220;
aud[31571]=16'he20d;
aud[31572]=16'he1fa;
aud[31573]=16'he1e8;
aud[31574]=16'he1d5;
aud[31575]=16'he1c2;
aud[31576]=16'he1af;
aud[31577]=16'he19c;
aud[31578]=16'he189;
aud[31579]=16'he176;
aud[31580]=16'he163;
aud[31581]=16'he151;
aud[31582]=16'he13e;
aud[31583]=16'he12b;
aud[31584]=16'he118;
aud[31585]=16'he105;
aud[31586]=16'he0f3;
aud[31587]=16'he0e0;
aud[31588]=16'he0cd;
aud[31589]=16'he0ba;
aud[31590]=16'he0a8;
aud[31591]=16'he095;
aud[31592]=16'he082;
aud[31593]=16'he070;
aud[31594]=16'he05d;
aud[31595]=16'he04a;
aud[31596]=16'he038;
aud[31597]=16'he025;
aud[31598]=16'he013;
aud[31599]=16'he000;
aud[31600]=16'hdfed;
aud[31601]=16'hdfdb;
aud[31602]=16'hdfc8;
aud[31603]=16'hdfb6;
aud[31604]=16'hdfa3;
aud[31605]=16'hdf91;
aud[31606]=16'hdf7e;
aud[31607]=16'hdf6c;
aud[31608]=16'hdf59;
aud[31609]=16'hdf47;
aud[31610]=16'hdf35;
aud[31611]=16'hdf22;
aud[31612]=16'hdf10;
aud[31613]=16'hdefd;
aud[31614]=16'hdeeb;
aud[31615]=16'hded9;
aud[31616]=16'hdec6;
aud[31617]=16'hdeb4;
aud[31618]=16'hdea2;
aud[31619]=16'hde8f;
aud[31620]=16'hde7d;
aud[31621]=16'hde6b;
aud[31622]=16'hde59;
aud[31623]=16'hde46;
aud[31624]=16'hde34;
aud[31625]=16'hde22;
aud[31626]=16'hde10;
aud[31627]=16'hddfe;
aud[31628]=16'hddeb;
aud[31629]=16'hddd9;
aud[31630]=16'hddc7;
aud[31631]=16'hddb5;
aud[31632]=16'hdda3;
aud[31633]=16'hdd91;
aud[31634]=16'hdd7f;
aud[31635]=16'hdd6d;
aud[31636]=16'hdd5b;
aud[31637]=16'hdd49;
aud[31638]=16'hdd37;
aud[31639]=16'hdd25;
aud[31640]=16'hdd13;
aud[31641]=16'hdd01;
aud[31642]=16'hdcef;
aud[31643]=16'hdcdd;
aud[31644]=16'hdccb;
aud[31645]=16'hdcb9;
aud[31646]=16'hdca7;
aud[31647]=16'hdc95;
aud[31648]=16'hdc83;
aud[31649]=16'hdc72;
aud[31650]=16'hdc60;
aud[31651]=16'hdc4e;
aud[31652]=16'hdc3c;
aud[31653]=16'hdc2a;
aud[31654]=16'hdc19;
aud[31655]=16'hdc07;
aud[31656]=16'hdbf5;
aud[31657]=16'hdbe3;
aud[31658]=16'hdbd2;
aud[31659]=16'hdbc0;
aud[31660]=16'hdbae;
aud[31661]=16'hdb9d;
aud[31662]=16'hdb8b;
aud[31663]=16'hdb79;
aud[31664]=16'hdb68;
aud[31665]=16'hdb56;
aud[31666]=16'hdb45;
aud[31667]=16'hdb33;
aud[31668]=16'hdb22;
aud[31669]=16'hdb10;
aud[31670]=16'hdaff;
aud[31671]=16'hdaed;
aud[31672]=16'hdadc;
aud[31673]=16'hdaca;
aud[31674]=16'hdab9;
aud[31675]=16'hdaa7;
aud[31676]=16'hda96;
aud[31677]=16'hda84;
aud[31678]=16'hda73;
aud[31679]=16'hda62;
aud[31680]=16'hda50;
aud[31681]=16'hda3f;
aud[31682]=16'hda2e;
aud[31683]=16'hda1c;
aud[31684]=16'hda0b;
aud[31685]=16'hd9fa;
aud[31686]=16'hd9e9;
aud[31687]=16'hd9d7;
aud[31688]=16'hd9c6;
aud[31689]=16'hd9b5;
aud[31690]=16'hd9a4;
aud[31691]=16'hd993;
aud[31692]=16'hd982;
aud[31693]=16'hd970;
aud[31694]=16'hd95f;
aud[31695]=16'hd94e;
aud[31696]=16'hd93d;
aud[31697]=16'hd92c;
aud[31698]=16'hd91b;
aud[31699]=16'hd90a;
aud[31700]=16'hd8f9;
aud[31701]=16'hd8e8;
aud[31702]=16'hd8d7;
aud[31703]=16'hd8c6;
aud[31704]=16'hd8b5;
aud[31705]=16'hd8a4;
aud[31706]=16'hd893;
aud[31707]=16'hd882;
aud[31708]=16'hd872;
aud[31709]=16'hd861;
aud[31710]=16'hd850;
aud[31711]=16'hd83f;
aud[31712]=16'hd82e;
aud[31713]=16'hd81e;
aud[31714]=16'hd80d;
aud[31715]=16'hd7fc;
aud[31716]=16'hd7eb;
aud[31717]=16'hd7db;
aud[31718]=16'hd7ca;
aud[31719]=16'hd7b9;
aud[31720]=16'hd7a9;
aud[31721]=16'hd798;
aud[31722]=16'hd787;
aud[31723]=16'hd777;
aud[31724]=16'hd766;
aud[31725]=16'hd756;
aud[31726]=16'hd745;
aud[31727]=16'hd734;
aud[31728]=16'hd724;
aud[31729]=16'hd713;
aud[31730]=16'hd703;
aud[31731]=16'hd6f2;
aud[31732]=16'hd6e2;
aud[31733]=16'hd6d2;
aud[31734]=16'hd6c1;
aud[31735]=16'hd6b1;
aud[31736]=16'hd6a0;
aud[31737]=16'hd690;
aud[31738]=16'hd680;
aud[31739]=16'hd66f;
aud[31740]=16'hd65f;
aud[31741]=16'hd64f;
aud[31742]=16'hd63f;
aud[31743]=16'hd62e;
aud[31744]=16'hd61e;
aud[31745]=16'hd60e;
aud[31746]=16'hd5fe;
aud[31747]=16'hd5ee;
aud[31748]=16'hd5dd;
aud[31749]=16'hd5cd;
aud[31750]=16'hd5bd;
aud[31751]=16'hd5ad;
aud[31752]=16'hd59d;
aud[31753]=16'hd58d;
aud[31754]=16'hd57d;
aud[31755]=16'hd56d;
aud[31756]=16'hd55d;
aud[31757]=16'hd54d;
aud[31758]=16'hd53d;
aud[31759]=16'hd52d;
aud[31760]=16'hd51d;
aud[31761]=16'hd50d;
aud[31762]=16'hd4fd;
aud[31763]=16'hd4ed;
aud[31764]=16'hd4de;
aud[31765]=16'hd4ce;
aud[31766]=16'hd4be;
aud[31767]=16'hd4ae;
aud[31768]=16'hd49e;
aud[31769]=16'hd48f;
aud[31770]=16'hd47f;
aud[31771]=16'hd46f;
aud[31772]=16'hd45f;
aud[31773]=16'hd450;
aud[31774]=16'hd440;
aud[31775]=16'hd430;
aud[31776]=16'hd421;
aud[31777]=16'hd411;
aud[31778]=16'hd402;
aud[31779]=16'hd3f2;
aud[31780]=16'hd3e2;
aud[31781]=16'hd3d3;
aud[31782]=16'hd3c3;
aud[31783]=16'hd3b4;
aud[31784]=16'hd3a4;
aud[31785]=16'hd395;
aud[31786]=16'hd386;
aud[31787]=16'hd376;
aud[31788]=16'hd367;
aud[31789]=16'hd357;
aud[31790]=16'hd348;
aud[31791]=16'hd339;
aud[31792]=16'hd329;
aud[31793]=16'hd31a;
aud[31794]=16'hd30b;
aud[31795]=16'hd2fc;
aud[31796]=16'hd2ec;
aud[31797]=16'hd2dd;
aud[31798]=16'hd2ce;
aud[31799]=16'hd2bf;
aud[31800]=16'hd2b0;
aud[31801]=16'hd2a0;
aud[31802]=16'hd291;
aud[31803]=16'hd282;
aud[31804]=16'hd273;
aud[31805]=16'hd264;
aud[31806]=16'hd255;
aud[31807]=16'hd246;
aud[31808]=16'hd237;
aud[31809]=16'hd228;
aud[31810]=16'hd219;
aud[31811]=16'hd20a;
aud[31812]=16'hd1fb;
aud[31813]=16'hd1ec;
aud[31814]=16'hd1de;
aud[31815]=16'hd1cf;
aud[31816]=16'hd1c0;
aud[31817]=16'hd1b1;
aud[31818]=16'hd1a2;
aud[31819]=16'hd193;
aud[31820]=16'hd185;
aud[31821]=16'hd176;
aud[31822]=16'hd167;
aud[31823]=16'hd159;
aud[31824]=16'hd14a;
aud[31825]=16'hd13b;
aud[31826]=16'hd12d;
aud[31827]=16'hd11e;
aud[31828]=16'hd10f;
aud[31829]=16'hd101;
aud[31830]=16'hd0f2;
aud[31831]=16'hd0e4;
aud[31832]=16'hd0d5;
aud[31833]=16'hd0c7;
aud[31834]=16'hd0b8;
aud[31835]=16'hd0aa;
aud[31836]=16'hd09b;
aud[31837]=16'hd08d;
aud[31838]=16'hd07f;
aud[31839]=16'hd070;
aud[31840]=16'hd062;
aud[31841]=16'hd054;
aud[31842]=16'hd045;
aud[31843]=16'hd037;
aud[31844]=16'hd029;
aud[31845]=16'hd01b;
aud[31846]=16'hd00c;
aud[31847]=16'hcffe;
aud[31848]=16'hcff0;
aud[31849]=16'hcfe2;
aud[31850]=16'hcfd4;
aud[31851]=16'hcfc6;
aud[31852]=16'hcfb8;
aud[31853]=16'hcfa9;
aud[31854]=16'hcf9b;
aud[31855]=16'hcf8d;
aud[31856]=16'hcf7f;
aud[31857]=16'hcf71;
aud[31858]=16'hcf63;
aud[31859]=16'hcf56;
aud[31860]=16'hcf48;
aud[31861]=16'hcf3a;
aud[31862]=16'hcf2c;
aud[31863]=16'hcf1e;
aud[31864]=16'hcf10;
aud[31865]=16'hcf02;
aud[31866]=16'hcef5;
aud[31867]=16'hcee7;
aud[31868]=16'hced9;
aud[31869]=16'hcecb;
aud[31870]=16'hcebe;
aud[31871]=16'hceb0;
aud[31872]=16'hcea2;
aud[31873]=16'hce95;
aud[31874]=16'hce87;
aud[31875]=16'hce79;
aud[31876]=16'hce6c;
aud[31877]=16'hce5e;
aud[31878]=16'hce51;
aud[31879]=16'hce43;
aud[31880]=16'hce36;
aud[31881]=16'hce28;
aud[31882]=16'hce1b;
aud[31883]=16'hce0d;
aud[31884]=16'hce00;
aud[31885]=16'hcdf3;
aud[31886]=16'hcde5;
aud[31887]=16'hcdd8;
aud[31888]=16'hcdcb;
aud[31889]=16'hcdbd;
aud[31890]=16'hcdb0;
aud[31891]=16'hcda3;
aud[31892]=16'hcd96;
aud[31893]=16'hcd88;
aud[31894]=16'hcd7b;
aud[31895]=16'hcd6e;
aud[31896]=16'hcd61;
aud[31897]=16'hcd54;
aud[31898]=16'hcd47;
aud[31899]=16'hcd3a;
aud[31900]=16'hcd2d;
aud[31901]=16'hcd20;
aud[31902]=16'hcd13;
aud[31903]=16'hcd06;
aud[31904]=16'hccf9;
aud[31905]=16'hccec;
aud[31906]=16'hccdf;
aud[31907]=16'hccd2;
aud[31908]=16'hccc5;
aud[31909]=16'hccb8;
aud[31910]=16'hccab;
aud[31911]=16'hcc9f;
aud[31912]=16'hcc92;
aud[31913]=16'hcc85;
aud[31914]=16'hcc78;
aud[31915]=16'hcc6c;
aud[31916]=16'hcc5f;
aud[31917]=16'hcc52;
aud[31918]=16'hcc46;
aud[31919]=16'hcc39;
aud[31920]=16'hcc2c;
aud[31921]=16'hcc20;
aud[31922]=16'hcc13;
aud[31923]=16'hcc07;
aud[31924]=16'hcbfa;
aud[31925]=16'hcbee;
aud[31926]=16'hcbe1;
aud[31927]=16'hcbd5;
aud[31928]=16'hcbc9;
aud[31929]=16'hcbbc;
aud[31930]=16'hcbb0;
aud[31931]=16'hcba3;
aud[31932]=16'hcb97;
aud[31933]=16'hcb8b;
aud[31934]=16'hcb7f;
aud[31935]=16'hcb72;
aud[31936]=16'hcb66;
aud[31937]=16'hcb5a;
aud[31938]=16'hcb4e;
aud[31939]=16'hcb42;
aud[31940]=16'hcb35;
aud[31941]=16'hcb29;
aud[31942]=16'hcb1d;
aud[31943]=16'hcb11;
aud[31944]=16'hcb05;
aud[31945]=16'hcaf9;
aud[31946]=16'hcaed;
aud[31947]=16'hcae1;
aud[31948]=16'hcad5;
aud[31949]=16'hcac9;
aud[31950]=16'hcabd;
aud[31951]=16'hcab1;
aud[31952]=16'hcaa6;
aud[31953]=16'hca9a;
aud[31954]=16'hca8e;
aud[31955]=16'hca82;
aud[31956]=16'hca76;
aud[31957]=16'hca6b;
aud[31958]=16'hca5f;
aud[31959]=16'hca53;
aud[31960]=16'hca48;
aud[31961]=16'hca3c;
aud[31962]=16'hca30;
aud[31963]=16'hca25;
aud[31964]=16'hca19;
aud[31965]=16'hca0e;
aud[31966]=16'hca02;
aud[31967]=16'hc9f7;
aud[31968]=16'hc9eb;
aud[31969]=16'hc9e0;
aud[31970]=16'hc9d4;
aud[31971]=16'hc9c9;
aud[31972]=16'hc9bd;
aud[31973]=16'hc9b2;
aud[31974]=16'hc9a7;
aud[31975]=16'hc99b;
aud[31976]=16'hc990;
aud[31977]=16'hc985;
aud[31978]=16'hc97a;
aud[31979]=16'hc96e;
aud[31980]=16'hc963;
aud[31981]=16'hc958;
aud[31982]=16'hc94d;
aud[31983]=16'hc942;
aud[31984]=16'hc937;
aud[31985]=16'hc92c;
aud[31986]=16'hc920;
aud[31987]=16'hc915;
aud[31988]=16'hc90a;
aud[31989]=16'hc8ff;
aud[31990]=16'hc8f5;
aud[31991]=16'hc8ea;
aud[31992]=16'hc8df;
aud[31993]=16'hc8d4;
aud[31994]=16'hc8c9;
aud[31995]=16'hc8be;
aud[31996]=16'hc8b3;
aud[31997]=16'hc8a9;
aud[31998]=16'hc89e;
aud[31999]=16'hc893;
aud[32000]=16'hc888;
aud[32001]=16'hc87e;
aud[32002]=16'hc873;
aud[32003]=16'hc868;
aud[32004]=16'hc85e;
aud[32005]=16'hc853;
aud[32006]=16'hc849;
aud[32007]=16'hc83e;
aud[32008]=16'hc834;
aud[32009]=16'hc829;
aud[32010]=16'hc81f;
aud[32011]=16'hc814;
aud[32012]=16'hc80a;
aud[32013]=16'hc7ff;
aud[32014]=16'hc7f5;
aud[32015]=16'hc7eb;
aud[32016]=16'hc7e0;
aud[32017]=16'hc7d6;
aud[32018]=16'hc7cc;
aud[32019]=16'hc7c1;
aud[32020]=16'hc7b7;
aud[32021]=16'hc7ad;
aud[32022]=16'hc7a3;
aud[32023]=16'hc799;
aud[32024]=16'hc78f;
aud[32025]=16'hc785;
aud[32026]=16'hc77a;
aud[32027]=16'hc770;
aud[32028]=16'hc766;
aud[32029]=16'hc75c;
aud[32030]=16'hc752;
aud[32031]=16'hc748;
aud[32032]=16'hc73f;
aud[32033]=16'hc735;
aud[32034]=16'hc72b;
aud[32035]=16'hc721;
aud[32036]=16'hc717;
aud[32037]=16'hc70d;
aud[32038]=16'hc703;
aud[32039]=16'hc6fa;
aud[32040]=16'hc6f0;
aud[32041]=16'hc6e6;
aud[32042]=16'hc6dd;
aud[32043]=16'hc6d3;
aud[32044]=16'hc6c9;
aud[32045]=16'hc6c0;
aud[32046]=16'hc6b6;
aud[32047]=16'hc6ad;
aud[32048]=16'hc6a3;
aud[32049]=16'hc69a;
aud[32050]=16'hc690;
aud[32051]=16'hc687;
aud[32052]=16'hc67d;
aud[32053]=16'hc674;
aud[32054]=16'hc66b;
aud[32055]=16'hc661;
aud[32056]=16'hc658;
aud[32057]=16'hc64f;
aud[32058]=16'hc645;
aud[32059]=16'hc63c;
aud[32060]=16'hc633;
aud[32061]=16'hc62a;
aud[32062]=16'hc620;
aud[32063]=16'hc617;
aud[32064]=16'hc60e;
aud[32065]=16'hc605;
aud[32066]=16'hc5fc;
aud[32067]=16'hc5f3;
aud[32068]=16'hc5ea;
aud[32069]=16'hc5e1;
aud[32070]=16'hc5d8;
aud[32071]=16'hc5cf;
aud[32072]=16'hc5c6;
aud[32073]=16'hc5bd;
aud[32074]=16'hc5b4;
aud[32075]=16'hc5ac;
aud[32076]=16'hc5a3;
aud[32077]=16'hc59a;
aud[32078]=16'hc591;
aud[32079]=16'hc588;
aud[32080]=16'hc580;
aud[32081]=16'hc577;
aud[32082]=16'hc56e;
aud[32083]=16'hc566;
aud[32084]=16'hc55d;
aud[32085]=16'hc555;
aud[32086]=16'hc54c;
aud[32087]=16'hc544;
aud[32088]=16'hc53b;
aud[32089]=16'hc533;
aud[32090]=16'hc52a;
aud[32091]=16'hc522;
aud[32092]=16'hc519;
aud[32093]=16'hc511;
aud[32094]=16'hc509;
aud[32095]=16'hc500;
aud[32096]=16'hc4f8;
aud[32097]=16'hc4f0;
aud[32098]=16'hc4e7;
aud[32099]=16'hc4df;
aud[32100]=16'hc4d7;
aud[32101]=16'hc4cf;
aud[32102]=16'hc4c7;
aud[32103]=16'hc4bf;
aud[32104]=16'hc4b6;
aud[32105]=16'hc4ae;
aud[32106]=16'hc4a6;
aud[32107]=16'hc49e;
aud[32108]=16'hc496;
aud[32109]=16'hc48e;
aud[32110]=16'hc486;
aud[32111]=16'hc47f;
aud[32112]=16'hc477;
aud[32113]=16'hc46f;
aud[32114]=16'hc467;
aud[32115]=16'hc45f;
aud[32116]=16'hc457;
aud[32117]=16'hc450;
aud[32118]=16'hc448;
aud[32119]=16'hc440;
aud[32120]=16'hc439;
aud[32121]=16'hc431;
aud[32122]=16'hc429;
aud[32123]=16'hc422;
aud[32124]=16'hc41a;
aud[32125]=16'hc413;
aud[32126]=16'hc40b;
aud[32127]=16'hc404;
aud[32128]=16'hc3fc;
aud[32129]=16'hc3f5;
aud[32130]=16'hc3ed;
aud[32131]=16'hc3e6;
aud[32132]=16'hc3df;
aud[32133]=16'hc3d7;
aud[32134]=16'hc3d0;
aud[32135]=16'hc3c9;
aud[32136]=16'hc3c1;
aud[32137]=16'hc3ba;
aud[32138]=16'hc3b3;
aud[32139]=16'hc3ac;
aud[32140]=16'hc3a5;
aud[32141]=16'hc39d;
aud[32142]=16'hc396;
aud[32143]=16'hc38f;
aud[32144]=16'hc388;
aud[32145]=16'hc381;
aud[32146]=16'hc37a;
aud[32147]=16'hc373;
aud[32148]=16'hc36c;
aud[32149]=16'hc365;
aud[32150]=16'hc35f;
aud[32151]=16'hc358;
aud[32152]=16'hc351;
aud[32153]=16'hc34a;
aud[32154]=16'hc343;
aud[32155]=16'hc33d;
aud[32156]=16'hc336;
aud[32157]=16'hc32f;
aud[32158]=16'hc329;
aud[32159]=16'hc322;
aud[32160]=16'hc31b;
aud[32161]=16'hc315;
aud[32162]=16'hc30e;
aud[32163]=16'hc308;
aud[32164]=16'hc301;
aud[32165]=16'hc2fb;
aud[32166]=16'hc2f4;
aud[32167]=16'hc2ee;
aud[32168]=16'hc2e7;
aud[32169]=16'hc2e1;
aud[32170]=16'hc2db;
aud[32171]=16'hc2d4;
aud[32172]=16'hc2ce;
aud[32173]=16'hc2c8;
aud[32174]=16'hc2c1;
aud[32175]=16'hc2bb;
aud[32176]=16'hc2b5;
aud[32177]=16'hc2af;
aud[32178]=16'hc2a9;
aud[32179]=16'hc2a3;
aud[32180]=16'hc29d;
aud[32181]=16'hc297;
aud[32182]=16'hc291;
aud[32183]=16'hc28b;
aud[32184]=16'hc285;
aud[32185]=16'hc27f;
aud[32186]=16'hc279;
aud[32187]=16'hc273;
aud[32188]=16'hc26d;
aud[32189]=16'hc267;
aud[32190]=16'hc261;
aud[32191]=16'hc25c;
aud[32192]=16'hc256;
aud[32193]=16'hc250;
aud[32194]=16'hc24a;
aud[32195]=16'hc245;
aud[32196]=16'hc23f;
aud[32197]=16'hc239;
aud[32198]=16'hc234;
aud[32199]=16'hc22e;
aud[32200]=16'hc229;
aud[32201]=16'hc223;
aud[32202]=16'hc21e;
aud[32203]=16'hc218;
aud[32204]=16'hc213;
aud[32205]=16'hc20d;
aud[32206]=16'hc208;
aud[32207]=16'hc203;
aud[32208]=16'hc1fd;
aud[32209]=16'hc1f8;
aud[32210]=16'hc1f3;
aud[32211]=16'hc1ee;
aud[32212]=16'hc1e8;
aud[32213]=16'hc1e3;
aud[32214]=16'hc1de;
aud[32215]=16'hc1d9;
aud[32216]=16'hc1d4;
aud[32217]=16'hc1cf;
aud[32218]=16'hc1ca;
aud[32219]=16'hc1c5;
aud[32220]=16'hc1c0;
aud[32221]=16'hc1bb;
aud[32222]=16'hc1b6;
aud[32223]=16'hc1b1;
aud[32224]=16'hc1ac;
aud[32225]=16'hc1a7;
aud[32226]=16'hc1a2;
aud[32227]=16'hc19e;
aud[32228]=16'hc199;
aud[32229]=16'hc194;
aud[32230]=16'hc18f;
aud[32231]=16'hc18b;
aud[32232]=16'hc186;
aud[32233]=16'hc181;
aud[32234]=16'hc17d;
aud[32235]=16'hc178;
aud[32236]=16'hc174;
aud[32237]=16'hc16f;
aud[32238]=16'hc16b;
aud[32239]=16'hc166;
aud[32240]=16'hc162;
aud[32241]=16'hc15d;
aud[32242]=16'hc159;
aud[32243]=16'hc154;
aud[32244]=16'hc150;
aud[32245]=16'hc14c;
aud[32246]=16'hc147;
aud[32247]=16'hc143;
aud[32248]=16'hc13f;
aud[32249]=16'hc13b;
aud[32250]=16'hc137;
aud[32251]=16'hc133;
aud[32252]=16'hc12e;
aud[32253]=16'hc12a;
aud[32254]=16'hc126;
aud[32255]=16'hc122;
aud[32256]=16'hc11e;
aud[32257]=16'hc11a;
aud[32258]=16'hc116;
aud[32259]=16'hc112;
aud[32260]=16'hc10e;
aud[32261]=16'hc10b;
aud[32262]=16'hc107;
aud[32263]=16'hc103;
aud[32264]=16'hc0ff;
aud[32265]=16'hc0fb;
aud[32266]=16'hc0f8;
aud[32267]=16'hc0f4;
aud[32268]=16'hc0f0;
aud[32269]=16'hc0ed;
aud[32270]=16'hc0e9;
aud[32271]=16'hc0e5;
aud[32272]=16'hc0e2;
aud[32273]=16'hc0de;
aud[32274]=16'hc0db;
aud[32275]=16'hc0d7;
aud[32276]=16'hc0d4;
aud[32277]=16'hc0d0;
aud[32278]=16'hc0cd;
aud[32279]=16'hc0ca;
aud[32280]=16'hc0c6;
aud[32281]=16'hc0c3;
aud[32282]=16'hc0c0;
aud[32283]=16'hc0bd;
aud[32284]=16'hc0b9;
aud[32285]=16'hc0b6;
aud[32286]=16'hc0b3;
aud[32287]=16'hc0b0;
aud[32288]=16'hc0ad;
aud[32289]=16'hc0aa;
aud[32290]=16'hc0a6;
aud[32291]=16'hc0a3;
aud[32292]=16'hc0a0;
aud[32293]=16'hc09d;
aud[32294]=16'hc09b;
aud[32295]=16'hc098;
aud[32296]=16'hc095;
aud[32297]=16'hc092;
aud[32298]=16'hc08f;
aud[32299]=16'hc08c;
aud[32300]=16'hc089;
aud[32301]=16'hc087;
aud[32302]=16'hc084;
aud[32303]=16'hc081;
aud[32304]=16'hc07f;
aud[32305]=16'hc07c;
aud[32306]=16'hc079;
aud[32307]=16'hc077;
aud[32308]=16'hc074;
aud[32309]=16'hc072;
aud[32310]=16'hc06f;
aud[32311]=16'hc06d;
aud[32312]=16'hc06a;
aud[32313]=16'hc068;
aud[32314]=16'hc065;
aud[32315]=16'hc063;
aud[32316]=16'hc061;
aud[32317]=16'hc05e;
aud[32318]=16'hc05c;
aud[32319]=16'hc05a;
aud[32320]=16'hc058;
aud[32321]=16'hc055;
aud[32322]=16'hc053;
aud[32323]=16'hc051;
aud[32324]=16'hc04f;
aud[32325]=16'hc04d;
aud[32326]=16'hc04b;
aud[32327]=16'hc049;
aud[32328]=16'hc047;
aud[32329]=16'hc045;
aud[32330]=16'hc043;
aud[32331]=16'hc041;
aud[32332]=16'hc03f;
aud[32333]=16'hc03d;
aud[32334]=16'hc03b;
aud[32335]=16'hc039;
aud[32336]=16'hc038;
aud[32337]=16'hc036;
aud[32338]=16'hc034;
aud[32339]=16'hc033;
aud[32340]=16'hc031;
aud[32341]=16'hc02f;
aud[32342]=16'hc02e;
aud[32343]=16'hc02c;
aud[32344]=16'hc02a;
aud[32345]=16'hc029;
aud[32346]=16'hc027;
aud[32347]=16'hc026;
aud[32348]=16'hc024;
aud[32349]=16'hc023;
aud[32350]=16'hc022;
aud[32351]=16'hc020;
aud[32352]=16'hc01f;
aud[32353]=16'hc01e;
aud[32354]=16'hc01c;
aud[32355]=16'hc01b;
aud[32356]=16'hc01a;
aud[32357]=16'hc019;
aud[32358]=16'hc018;
aud[32359]=16'hc016;
aud[32360]=16'hc015;
aud[32361]=16'hc014;
aud[32362]=16'hc013;
aud[32363]=16'hc012;
aud[32364]=16'hc011;
aud[32365]=16'hc010;
aud[32366]=16'hc00f;
aud[32367]=16'hc00e;
aud[32368]=16'hc00d;
aud[32369]=16'hc00d;
aud[32370]=16'hc00c;
aud[32371]=16'hc00b;
aud[32372]=16'hc00a;
aud[32373]=16'hc009;
aud[32374]=16'hc009;
aud[32375]=16'hc008;
aud[32376]=16'hc007;
aud[32377]=16'hc007;
aud[32378]=16'hc006;
aud[32379]=16'hc006;
aud[32380]=16'hc005;
aud[32381]=16'hc005;
aud[32382]=16'hc004;
aud[32383]=16'hc004;
aud[32384]=16'hc003;
aud[32385]=16'hc003;
aud[32386]=16'hc002;
aud[32387]=16'hc002;
aud[32388]=16'hc002;
aud[32389]=16'hc001;
aud[32390]=16'hc001;
aud[32391]=16'hc001;
aud[32392]=16'hc001;
aud[32393]=16'hc001;
aud[32394]=16'hc000;
aud[32395]=16'hc000;
aud[32396]=16'hc000;
aud[32397]=16'hc000;
aud[32398]=16'hc000;
aud[32399]=16'hc000;
aud[32400]=16'hc000;
aud[32401]=16'hc000;
aud[32402]=16'hc000;
aud[32403]=16'hc000;
aud[32404]=16'hc000;
aud[32405]=16'hc001;
aud[32406]=16'hc001;
aud[32407]=16'hc001;
aud[32408]=16'hc001;
aud[32409]=16'hc001;
aud[32410]=16'hc002;
aud[32411]=16'hc002;
aud[32412]=16'hc002;
aud[32413]=16'hc003;
aud[32414]=16'hc003;
aud[32415]=16'hc004;
aud[32416]=16'hc004;
aud[32417]=16'hc005;
aud[32418]=16'hc005;
aud[32419]=16'hc006;
aud[32420]=16'hc006;
aud[32421]=16'hc007;
aud[32422]=16'hc007;
aud[32423]=16'hc008;
aud[32424]=16'hc009;
aud[32425]=16'hc009;
aud[32426]=16'hc00a;
aud[32427]=16'hc00b;
aud[32428]=16'hc00c;
aud[32429]=16'hc00d;
aud[32430]=16'hc00d;
aud[32431]=16'hc00e;
aud[32432]=16'hc00f;
aud[32433]=16'hc010;
aud[32434]=16'hc011;
aud[32435]=16'hc012;
aud[32436]=16'hc013;
aud[32437]=16'hc014;
aud[32438]=16'hc015;
aud[32439]=16'hc016;
aud[32440]=16'hc018;
aud[32441]=16'hc019;
aud[32442]=16'hc01a;
aud[32443]=16'hc01b;
aud[32444]=16'hc01c;
aud[32445]=16'hc01e;
aud[32446]=16'hc01f;
aud[32447]=16'hc020;
aud[32448]=16'hc022;
aud[32449]=16'hc023;
aud[32450]=16'hc024;
aud[32451]=16'hc026;
aud[32452]=16'hc027;
aud[32453]=16'hc029;
aud[32454]=16'hc02a;
aud[32455]=16'hc02c;
aud[32456]=16'hc02e;
aud[32457]=16'hc02f;
aud[32458]=16'hc031;
aud[32459]=16'hc033;
aud[32460]=16'hc034;
aud[32461]=16'hc036;
aud[32462]=16'hc038;
aud[32463]=16'hc039;
aud[32464]=16'hc03b;
aud[32465]=16'hc03d;
aud[32466]=16'hc03f;
aud[32467]=16'hc041;
aud[32468]=16'hc043;
aud[32469]=16'hc045;
aud[32470]=16'hc047;
aud[32471]=16'hc049;
aud[32472]=16'hc04b;
aud[32473]=16'hc04d;
aud[32474]=16'hc04f;
aud[32475]=16'hc051;
aud[32476]=16'hc053;
aud[32477]=16'hc055;
aud[32478]=16'hc058;
aud[32479]=16'hc05a;
aud[32480]=16'hc05c;
aud[32481]=16'hc05e;
aud[32482]=16'hc061;
aud[32483]=16'hc063;
aud[32484]=16'hc065;
aud[32485]=16'hc068;
aud[32486]=16'hc06a;
aud[32487]=16'hc06d;
aud[32488]=16'hc06f;
aud[32489]=16'hc072;
aud[32490]=16'hc074;
aud[32491]=16'hc077;
aud[32492]=16'hc079;
aud[32493]=16'hc07c;
aud[32494]=16'hc07f;
aud[32495]=16'hc081;
aud[32496]=16'hc084;
aud[32497]=16'hc087;
aud[32498]=16'hc089;
aud[32499]=16'hc08c;
aud[32500]=16'hc08f;
aud[32501]=16'hc092;
aud[32502]=16'hc095;
aud[32503]=16'hc098;
aud[32504]=16'hc09b;
aud[32505]=16'hc09d;
aud[32506]=16'hc0a0;
aud[32507]=16'hc0a3;
aud[32508]=16'hc0a6;
aud[32509]=16'hc0aa;
aud[32510]=16'hc0ad;
aud[32511]=16'hc0b0;
aud[32512]=16'hc0b3;
aud[32513]=16'hc0b6;
aud[32514]=16'hc0b9;
aud[32515]=16'hc0bd;
aud[32516]=16'hc0c0;
aud[32517]=16'hc0c3;
aud[32518]=16'hc0c6;
aud[32519]=16'hc0ca;
aud[32520]=16'hc0cd;
aud[32521]=16'hc0d0;
aud[32522]=16'hc0d4;
aud[32523]=16'hc0d7;
aud[32524]=16'hc0db;
aud[32525]=16'hc0de;
aud[32526]=16'hc0e2;
aud[32527]=16'hc0e5;
aud[32528]=16'hc0e9;
aud[32529]=16'hc0ed;
aud[32530]=16'hc0f0;
aud[32531]=16'hc0f4;
aud[32532]=16'hc0f8;
aud[32533]=16'hc0fb;
aud[32534]=16'hc0ff;
aud[32535]=16'hc103;
aud[32536]=16'hc107;
aud[32537]=16'hc10b;
aud[32538]=16'hc10e;
aud[32539]=16'hc112;
aud[32540]=16'hc116;
aud[32541]=16'hc11a;
aud[32542]=16'hc11e;
aud[32543]=16'hc122;
aud[32544]=16'hc126;
aud[32545]=16'hc12a;
aud[32546]=16'hc12e;
aud[32547]=16'hc133;
aud[32548]=16'hc137;
aud[32549]=16'hc13b;
aud[32550]=16'hc13f;
aud[32551]=16'hc143;
aud[32552]=16'hc147;
aud[32553]=16'hc14c;
aud[32554]=16'hc150;
aud[32555]=16'hc154;
aud[32556]=16'hc159;
aud[32557]=16'hc15d;
aud[32558]=16'hc162;
aud[32559]=16'hc166;
aud[32560]=16'hc16b;
aud[32561]=16'hc16f;
aud[32562]=16'hc174;
aud[32563]=16'hc178;
aud[32564]=16'hc17d;
aud[32565]=16'hc181;
aud[32566]=16'hc186;
aud[32567]=16'hc18b;
aud[32568]=16'hc18f;
aud[32569]=16'hc194;
aud[32570]=16'hc199;
aud[32571]=16'hc19e;
aud[32572]=16'hc1a2;
aud[32573]=16'hc1a7;
aud[32574]=16'hc1ac;
aud[32575]=16'hc1b1;
aud[32576]=16'hc1b6;
aud[32577]=16'hc1bb;
aud[32578]=16'hc1c0;
aud[32579]=16'hc1c5;
aud[32580]=16'hc1ca;
aud[32581]=16'hc1cf;
aud[32582]=16'hc1d4;
aud[32583]=16'hc1d9;
aud[32584]=16'hc1de;
aud[32585]=16'hc1e3;
aud[32586]=16'hc1e8;
aud[32587]=16'hc1ee;
aud[32588]=16'hc1f3;
aud[32589]=16'hc1f8;
aud[32590]=16'hc1fd;
aud[32591]=16'hc203;
aud[32592]=16'hc208;
aud[32593]=16'hc20d;
aud[32594]=16'hc213;
aud[32595]=16'hc218;
aud[32596]=16'hc21e;
aud[32597]=16'hc223;
aud[32598]=16'hc229;
aud[32599]=16'hc22e;
aud[32600]=16'hc234;
aud[32601]=16'hc239;
aud[32602]=16'hc23f;
aud[32603]=16'hc245;
aud[32604]=16'hc24a;
aud[32605]=16'hc250;
aud[32606]=16'hc256;
aud[32607]=16'hc25c;
aud[32608]=16'hc261;
aud[32609]=16'hc267;
aud[32610]=16'hc26d;
aud[32611]=16'hc273;
aud[32612]=16'hc279;
aud[32613]=16'hc27f;
aud[32614]=16'hc285;
aud[32615]=16'hc28b;
aud[32616]=16'hc291;
aud[32617]=16'hc297;
aud[32618]=16'hc29d;
aud[32619]=16'hc2a3;
aud[32620]=16'hc2a9;
aud[32621]=16'hc2af;
aud[32622]=16'hc2b5;
aud[32623]=16'hc2bb;
aud[32624]=16'hc2c1;
aud[32625]=16'hc2c8;
aud[32626]=16'hc2ce;
aud[32627]=16'hc2d4;
aud[32628]=16'hc2db;
aud[32629]=16'hc2e1;
aud[32630]=16'hc2e7;
aud[32631]=16'hc2ee;
aud[32632]=16'hc2f4;
aud[32633]=16'hc2fb;
aud[32634]=16'hc301;
aud[32635]=16'hc308;
aud[32636]=16'hc30e;
aud[32637]=16'hc315;
aud[32638]=16'hc31b;
aud[32639]=16'hc322;
aud[32640]=16'hc329;
aud[32641]=16'hc32f;
aud[32642]=16'hc336;
aud[32643]=16'hc33d;
aud[32644]=16'hc343;
aud[32645]=16'hc34a;
aud[32646]=16'hc351;
aud[32647]=16'hc358;
aud[32648]=16'hc35f;
aud[32649]=16'hc365;
aud[32650]=16'hc36c;
aud[32651]=16'hc373;
aud[32652]=16'hc37a;
aud[32653]=16'hc381;
aud[32654]=16'hc388;
aud[32655]=16'hc38f;
aud[32656]=16'hc396;
aud[32657]=16'hc39d;
aud[32658]=16'hc3a5;
aud[32659]=16'hc3ac;
aud[32660]=16'hc3b3;
aud[32661]=16'hc3ba;
aud[32662]=16'hc3c1;
aud[32663]=16'hc3c9;
aud[32664]=16'hc3d0;
aud[32665]=16'hc3d7;
aud[32666]=16'hc3df;
aud[32667]=16'hc3e6;
aud[32668]=16'hc3ed;
aud[32669]=16'hc3f5;
aud[32670]=16'hc3fc;
aud[32671]=16'hc404;
aud[32672]=16'hc40b;
aud[32673]=16'hc413;
aud[32674]=16'hc41a;
aud[32675]=16'hc422;
aud[32676]=16'hc429;
aud[32677]=16'hc431;
aud[32678]=16'hc439;
aud[32679]=16'hc440;
aud[32680]=16'hc448;
aud[32681]=16'hc450;
aud[32682]=16'hc457;
aud[32683]=16'hc45f;
aud[32684]=16'hc467;
aud[32685]=16'hc46f;
aud[32686]=16'hc477;
aud[32687]=16'hc47f;
aud[32688]=16'hc486;
aud[32689]=16'hc48e;
aud[32690]=16'hc496;
aud[32691]=16'hc49e;
aud[32692]=16'hc4a6;
aud[32693]=16'hc4ae;
aud[32694]=16'hc4b6;
aud[32695]=16'hc4bf;
aud[32696]=16'hc4c7;
aud[32697]=16'hc4cf;
aud[32698]=16'hc4d7;
aud[32699]=16'hc4df;
aud[32700]=16'hc4e7;
aud[32701]=16'hc4f0;
aud[32702]=16'hc4f8;
aud[32703]=16'hc500;
aud[32704]=16'hc509;
aud[32705]=16'hc511;
aud[32706]=16'hc519;
aud[32707]=16'hc522;
aud[32708]=16'hc52a;
aud[32709]=16'hc533;
aud[32710]=16'hc53b;
aud[32711]=16'hc544;
aud[32712]=16'hc54c;
aud[32713]=16'hc555;
aud[32714]=16'hc55d;
aud[32715]=16'hc566;
aud[32716]=16'hc56e;
aud[32717]=16'hc577;
aud[32718]=16'hc580;
aud[32719]=16'hc588;
aud[32720]=16'hc591;
aud[32721]=16'hc59a;
aud[32722]=16'hc5a3;
aud[32723]=16'hc5ac;
aud[32724]=16'hc5b4;
aud[32725]=16'hc5bd;
aud[32726]=16'hc5c6;
aud[32727]=16'hc5cf;
aud[32728]=16'hc5d8;
aud[32729]=16'hc5e1;
aud[32730]=16'hc5ea;
aud[32731]=16'hc5f3;
aud[32732]=16'hc5fc;
aud[32733]=16'hc605;
aud[32734]=16'hc60e;
aud[32735]=16'hc617;
aud[32736]=16'hc620;
aud[32737]=16'hc62a;
aud[32738]=16'hc633;
aud[32739]=16'hc63c;
aud[32740]=16'hc645;
aud[32741]=16'hc64f;
aud[32742]=16'hc658;
aud[32743]=16'hc661;
aud[32744]=16'hc66b;
aud[32745]=16'hc674;
aud[32746]=16'hc67d;
aud[32747]=16'hc687;
aud[32748]=16'hc690;
aud[32749]=16'hc69a;
aud[32750]=16'hc6a3;
aud[32751]=16'hc6ad;
aud[32752]=16'hc6b6;
aud[32753]=16'hc6c0;
aud[32754]=16'hc6c9;
aud[32755]=16'hc6d3;
aud[32756]=16'hc6dd;
aud[32757]=16'hc6e6;
aud[32758]=16'hc6f0;
aud[32759]=16'hc6fa;
aud[32760]=16'hc703;
aud[32761]=16'hc70d;
aud[32762]=16'hc717;
aud[32763]=16'hc721;
aud[32764]=16'hc72b;
aud[32765]=16'hc735;
aud[32766]=16'hc73f;
aud[32767]=16'hc748;
aud[32768]=16'hc752;
aud[32769]=16'hc75c;
aud[32770]=16'hc766;
aud[32771]=16'hc770;
aud[32772]=16'hc77a;
aud[32773]=16'hc785;
aud[32774]=16'hc78f;
aud[32775]=16'hc799;
aud[32776]=16'hc7a3;
aud[32777]=16'hc7ad;
aud[32778]=16'hc7b7;
aud[32779]=16'hc7c1;
aud[32780]=16'hc7cc;
aud[32781]=16'hc7d6;
aud[32782]=16'hc7e0;
aud[32783]=16'hc7eb;
aud[32784]=16'hc7f5;
aud[32785]=16'hc7ff;
aud[32786]=16'hc80a;
aud[32787]=16'hc814;
aud[32788]=16'hc81f;
aud[32789]=16'hc829;
aud[32790]=16'hc834;
aud[32791]=16'hc83e;
aud[32792]=16'hc849;
aud[32793]=16'hc853;
aud[32794]=16'hc85e;
aud[32795]=16'hc868;
aud[32796]=16'hc873;
aud[32797]=16'hc87e;
aud[32798]=16'hc888;
aud[32799]=16'hc893;
aud[32800]=16'hc89e;
aud[32801]=16'hc8a9;
aud[32802]=16'hc8b3;
aud[32803]=16'hc8be;
aud[32804]=16'hc8c9;
aud[32805]=16'hc8d4;
aud[32806]=16'hc8df;
aud[32807]=16'hc8ea;
aud[32808]=16'hc8f5;
aud[32809]=16'hc8ff;
aud[32810]=16'hc90a;
aud[32811]=16'hc915;
aud[32812]=16'hc920;
aud[32813]=16'hc92c;
aud[32814]=16'hc937;
aud[32815]=16'hc942;
aud[32816]=16'hc94d;
aud[32817]=16'hc958;
aud[32818]=16'hc963;
aud[32819]=16'hc96e;
aud[32820]=16'hc97a;
aud[32821]=16'hc985;
aud[32822]=16'hc990;
aud[32823]=16'hc99b;
aud[32824]=16'hc9a7;
aud[32825]=16'hc9b2;
aud[32826]=16'hc9bd;
aud[32827]=16'hc9c9;
aud[32828]=16'hc9d4;
aud[32829]=16'hc9e0;
aud[32830]=16'hc9eb;
aud[32831]=16'hc9f7;
aud[32832]=16'hca02;
aud[32833]=16'hca0e;
aud[32834]=16'hca19;
aud[32835]=16'hca25;
aud[32836]=16'hca30;
aud[32837]=16'hca3c;
aud[32838]=16'hca48;
aud[32839]=16'hca53;
aud[32840]=16'hca5f;
aud[32841]=16'hca6b;
aud[32842]=16'hca76;
aud[32843]=16'hca82;
aud[32844]=16'hca8e;
aud[32845]=16'hca9a;
aud[32846]=16'hcaa6;
aud[32847]=16'hcab1;
aud[32848]=16'hcabd;
aud[32849]=16'hcac9;
aud[32850]=16'hcad5;
aud[32851]=16'hcae1;
aud[32852]=16'hcaed;
aud[32853]=16'hcaf9;
aud[32854]=16'hcb05;
aud[32855]=16'hcb11;
aud[32856]=16'hcb1d;
aud[32857]=16'hcb29;
aud[32858]=16'hcb35;
aud[32859]=16'hcb42;
aud[32860]=16'hcb4e;
aud[32861]=16'hcb5a;
aud[32862]=16'hcb66;
aud[32863]=16'hcb72;
aud[32864]=16'hcb7f;
aud[32865]=16'hcb8b;
aud[32866]=16'hcb97;
aud[32867]=16'hcba3;
aud[32868]=16'hcbb0;
aud[32869]=16'hcbbc;
aud[32870]=16'hcbc9;
aud[32871]=16'hcbd5;
aud[32872]=16'hcbe1;
aud[32873]=16'hcbee;
aud[32874]=16'hcbfa;
aud[32875]=16'hcc07;
aud[32876]=16'hcc13;
aud[32877]=16'hcc20;
aud[32878]=16'hcc2c;
aud[32879]=16'hcc39;
aud[32880]=16'hcc46;
aud[32881]=16'hcc52;
aud[32882]=16'hcc5f;
aud[32883]=16'hcc6c;
aud[32884]=16'hcc78;
aud[32885]=16'hcc85;
aud[32886]=16'hcc92;
aud[32887]=16'hcc9f;
aud[32888]=16'hccab;
aud[32889]=16'hccb8;
aud[32890]=16'hccc5;
aud[32891]=16'hccd2;
aud[32892]=16'hccdf;
aud[32893]=16'hccec;
aud[32894]=16'hccf9;
aud[32895]=16'hcd06;
aud[32896]=16'hcd13;
aud[32897]=16'hcd20;
aud[32898]=16'hcd2d;
aud[32899]=16'hcd3a;
aud[32900]=16'hcd47;
aud[32901]=16'hcd54;
aud[32902]=16'hcd61;
aud[32903]=16'hcd6e;
aud[32904]=16'hcd7b;
aud[32905]=16'hcd88;
aud[32906]=16'hcd96;
aud[32907]=16'hcda3;
aud[32908]=16'hcdb0;
aud[32909]=16'hcdbd;
aud[32910]=16'hcdcb;
aud[32911]=16'hcdd8;
aud[32912]=16'hcde5;
aud[32913]=16'hcdf3;
aud[32914]=16'hce00;
aud[32915]=16'hce0d;
aud[32916]=16'hce1b;
aud[32917]=16'hce28;
aud[32918]=16'hce36;
aud[32919]=16'hce43;
aud[32920]=16'hce51;
aud[32921]=16'hce5e;
aud[32922]=16'hce6c;
aud[32923]=16'hce79;
aud[32924]=16'hce87;
aud[32925]=16'hce95;
aud[32926]=16'hcea2;
aud[32927]=16'hceb0;
aud[32928]=16'hcebe;
aud[32929]=16'hcecb;
aud[32930]=16'hced9;
aud[32931]=16'hcee7;
aud[32932]=16'hcef5;
aud[32933]=16'hcf02;
aud[32934]=16'hcf10;
aud[32935]=16'hcf1e;
aud[32936]=16'hcf2c;
aud[32937]=16'hcf3a;
aud[32938]=16'hcf48;
aud[32939]=16'hcf56;
aud[32940]=16'hcf63;
aud[32941]=16'hcf71;
aud[32942]=16'hcf7f;
aud[32943]=16'hcf8d;
aud[32944]=16'hcf9b;
aud[32945]=16'hcfa9;
aud[32946]=16'hcfb8;
aud[32947]=16'hcfc6;
aud[32948]=16'hcfd4;
aud[32949]=16'hcfe2;
aud[32950]=16'hcff0;
aud[32951]=16'hcffe;
aud[32952]=16'hd00c;
aud[32953]=16'hd01b;
aud[32954]=16'hd029;
aud[32955]=16'hd037;
aud[32956]=16'hd045;
aud[32957]=16'hd054;
aud[32958]=16'hd062;
aud[32959]=16'hd070;
aud[32960]=16'hd07f;
aud[32961]=16'hd08d;
aud[32962]=16'hd09b;
aud[32963]=16'hd0aa;
aud[32964]=16'hd0b8;
aud[32965]=16'hd0c7;
aud[32966]=16'hd0d5;
aud[32967]=16'hd0e4;
aud[32968]=16'hd0f2;
aud[32969]=16'hd101;
aud[32970]=16'hd10f;
aud[32971]=16'hd11e;
aud[32972]=16'hd12d;
aud[32973]=16'hd13b;
aud[32974]=16'hd14a;
aud[32975]=16'hd159;
aud[32976]=16'hd167;
aud[32977]=16'hd176;
aud[32978]=16'hd185;
aud[32979]=16'hd193;
aud[32980]=16'hd1a2;
aud[32981]=16'hd1b1;
aud[32982]=16'hd1c0;
aud[32983]=16'hd1cf;
aud[32984]=16'hd1de;
aud[32985]=16'hd1ec;
aud[32986]=16'hd1fb;
aud[32987]=16'hd20a;
aud[32988]=16'hd219;
aud[32989]=16'hd228;
aud[32990]=16'hd237;
aud[32991]=16'hd246;
aud[32992]=16'hd255;
aud[32993]=16'hd264;
aud[32994]=16'hd273;
aud[32995]=16'hd282;
aud[32996]=16'hd291;
aud[32997]=16'hd2a0;
aud[32998]=16'hd2b0;
aud[32999]=16'hd2bf;
aud[33000]=16'hd2ce;
aud[33001]=16'hd2dd;
aud[33002]=16'hd2ec;
aud[33003]=16'hd2fc;
aud[33004]=16'hd30b;
aud[33005]=16'hd31a;
aud[33006]=16'hd329;
aud[33007]=16'hd339;
aud[33008]=16'hd348;
aud[33009]=16'hd357;
aud[33010]=16'hd367;
aud[33011]=16'hd376;
aud[33012]=16'hd386;
aud[33013]=16'hd395;
aud[33014]=16'hd3a4;
aud[33015]=16'hd3b4;
aud[33016]=16'hd3c3;
aud[33017]=16'hd3d3;
aud[33018]=16'hd3e2;
aud[33019]=16'hd3f2;
aud[33020]=16'hd402;
aud[33021]=16'hd411;
aud[33022]=16'hd421;
aud[33023]=16'hd430;
aud[33024]=16'hd440;
aud[33025]=16'hd450;
aud[33026]=16'hd45f;
aud[33027]=16'hd46f;
aud[33028]=16'hd47f;
aud[33029]=16'hd48f;
aud[33030]=16'hd49e;
aud[33031]=16'hd4ae;
aud[33032]=16'hd4be;
aud[33033]=16'hd4ce;
aud[33034]=16'hd4de;
aud[33035]=16'hd4ed;
aud[33036]=16'hd4fd;
aud[33037]=16'hd50d;
aud[33038]=16'hd51d;
aud[33039]=16'hd52d;
aud[33040]=16'hd53d;
aud[33041]=16'hd54d;
aud[33042]=16'hd55d;
aud[33043]=16'hd56d;
aud[33044]=16'hd57d;
aud[33045]=16'hd58d;
aud[33046]=16'hd59d;
aud[33047]=16'hd5ad;
aud[33048]=16'hd5bd;
aud[33049]=16'hd5cd;
aud[33050]=16'hd5dd;
aud[33051]=16'hd5ee;
aud[33052]=16'hd5fe;
aud[33053]=16'hd60e;
aud[33054]=16'hd61e;
aud[33055]=16'hd62e;
aud[33056]=16'hd63f;
aud[33057]=16'hd64f;
aud[33058]=16'hd65f;
aud[33059]=16'hd66f;
aud[33060]=16'hd680;
aud[33061]=16'hd690;
aud[33062]=16'hd6a0;
aud[33063]=16'hd6b1;
aud[33064]=16'hd6c1;
aud[33065]=16'hd6d2;
aud[33066]=16'hd6e2;
aud[33067]=16'hd6f2;
aud[33068]=16'hd703;
aud[33069]=16'hd713;
aud[33070]=16'hd724;
aud[33071]=16'hd734;
aud[33072]=16'hd745;
aud[33073]=16'hd756;
aud[33074]=16'hd766;
aud[33075]=16'hd777;
aud[33076]=16'hd787;
aud[33077]=16'hd798;
aud[33078]=16'hd7a9;
aud[33079]=16'hd7b9;
aud[33080]=16'hd7ca;
aud[33081]=16'hd7db;
aud[33082]=16'hd7eb;
aud[33083]=16'hd7fc;
aud[33084]=16'hd80d;
aud[33085]=16'hd81e;
aud[33086]=16'hd82e;
aud[33087]=16'hd83f;
aud[33088]=16'hd850;
aud[33089]=16'hd861;
aud[33090]=16'hd872;
aud[33091]=16'hd882;
aud[33092]=16'hd893;
aud[33093]=16'hd8a4;
aud[33094]=16'hd8b5;
aud[33095]=16'hd8c6;
aud[33096]=16'hd8d7;
aud[33097]=16'hd8e8;
aud[33098]=16'hd8f9;
aud[33099]=16'hd90a;
aud[33100]=16'hd91b;
aud[33101]=16'hd92c;
aud[33102]=16'hd93d;
aud[33103]=16'hd94e;
aud[33104]=16'hd95f;
aud[33105]=16'hd970;
aud[33106]=16'hd982;
aud[33107]=16'hd993;
aud[33108]=16'hd9a4;
aud[33109]=16'hd9b5;
aud[33110]=16'hd9c6;
aud[33111]=16'hd9d7;
aud[33112]=16'hd9e9;
aud[33113]=16'hd9fa;
aud[33114]=16'hda0b;
aud[33115]=16'hda1c;
aud[33116]=16'hda2e;
aud[33117]=16'hda3f;
aud[33118]=16'hda50;
aud[33119]=16'hda62;
aud[33120]=16'hda73;
aud[33121]=16'hda84;
aud[33122]=16'hda96;
aud[33123]=16'hdaa7;
aud[33124]=16'hdab9;
aud[33125]=16'hdaca;
aud[33126]=16'hdadc;
aud[33127]=16'hdaed;
aud[33128]=16'hdaff;
aud[33129]=16'hdb10;
aud[33130]=16'hdb22;
aud[33131]=16'hdb33;
aud[33132]=16'hdb45;
aud[33133]=16'hdb56;
aud[33134]=16'hdb68;
aud[33135]=16'hdb79;
aud[33136]=16'hdb8b;
aud[33137]=16'hdb9d;
aud[33138]=16'hdbae;
aud[33139]=16'hdbc0;
aud[33140]=16'hdbd2;
aud[33141]=16'hdbe3;
aud[33142]=16'hdbf5;
aud[33143]=16'hdc07;
aud[33144]=16'hdc19;
aud[33145]=16'hdc2a;
aud[33146]=16'hdc3c;
aud[33147]=16'hdc4e;
aud[33148]=16'hdc60;
aud[33149]=16'hdc72;
aud[33150]=16'hdc83;
aud[33151]=16'hdc95;
aud[33152]=16'hdca7;
aud[33153]=16'hdcb9;
aud[33154]=16'hdccb;
aud[33155]=16'hdcdd;
aud[33156]=16'hdcef;
aud[33157]=16'hdd01;
aud[33158]=16'hdd13;
aud[33159]=16'hdd25;
aud[33160]=16'hdd37;
aud[33161]=16'hdd49;
aud[33162]=16'hdd5b;
aud[33163]=16'hdd6d;
aud[33164]=16'hdd7f;
aud[33165]=16'hdd91;
aud[33166]=16'hdda3;
aud[33167]=16'hddb5;
aud[33168]=16'hddc7;
aud[33169]=16'hddd9;
aud[33170]=16'hddeb;
aud[33171]=16'hddfe;
aud[33172]=16'hde10;
aud[33173]=16'hde22;
aud[33174]=16'hde34;
aud[33175]=16'hde46;
aud[33176]=16'hde59;
aud[33177]=16'hde6b;
aud[33178]=16'hde7d;
aud[33179]=16'hde8f;
aud[33180]=16'hdea2;
aud[33181]=16'hdeb4;
aud[33182]=16'hdec6;
aud[33183]=16'hded9;
aud[33184]=16'hdeeb;
aud[33185]=16'hdefd;
aud[33186]=16'hdf10;
aud[33187]=16'hdf22;
aud[33188]=16'hdf35;
aud[33189]=16'hdf47;
aud[33190]=16'hdf59;
aud[33191]=16'hdf6c;
aud[33192]=16'hdf7e;
aud[33193]=16'hdf91;
aud[33194]=16'hdfa3;
aud[33195]=16'hdfb6;
aud[33196]=16'hdfc8;
aud[33197]=16'hdfdb;
aud[33198]=16'hdfed;
aud[33199]=16'he000;
aud[33200]=16'he013;
aud[33201]=16'he025;
aud[33202]=16'he038;
aud[33203]=16'he04a;
aud[33204]=16'he05d;
aud[33205]=16'he070;
aud[33206]=16'he082;
aud[33207]=16'he095;
aud[33208]=16'he0a8;
aud[33209]=16'he0ba;
aud[33210]=16'he0cd;
aud[33211]=16'he0e0;
aud[33212]=16'he0f3;
aud[33213]=16'he105;
aud[33214]=16'he118;
aud[33215]=16'he12b;
aud[33216]=16'he13e;
aud[33217]=16'he151;
aud[33218]=16'he163;
aud[33219]=16'he176;
aud[33220]=16'he189;
aud[33221]=16'he19c;
aud[33222]=16'he1af;
aud[33223]=16'he1c2;
aud[33224]=16'he1d5;
aud[33225]=16'he1e8;
aud[33226]=16'he1fa;
aud[33227]=16'he20d;
aud[33228]=16'he220;
aud[33229]=16'he233;
aud[33230]=16'he246;
aud[33231]=16'he259;
aud[33232]=16'he26c;
aud[33233]=16'he27f;
aud[33234]=16'he292;
aud[33235]=16'he2a5;
aud[33236]=16'he2b9;
aud[33237]=16'he2cc;
aud[33238]=16'he2df;
aud[33239]=16'he2f2;
aud[33240]=16'he305;
aud[33241]=16'he318;
aud[33242]=16'he32b;
aud[33243]=16'he33e;
aud[33244]=16'he352;
aud[33245]=16'he365;
aud[33246]=16'he378;
aud[33247]=16'he38b;
aud[33248]=16'he39e;
aud[33249]=16'he3b2;
aud[33250]=16'he3c5;
aud[33251]=16'he3d8;
aud[33252]=16'he3eb;
aud[33253]=16'he3ff;
aud[33254]=16'he412;
aud[33255]=16'he425;
aud[33256]=16'he438;
aud[33257]=16'he44c;
aud[33258]=16'he45f;
aud[33259]=16'he473;
aud[33260]=16'he486;
aud[33261]=16'he499;
aud[33262]=16'he4ad;
aud[33263]=16'he4c0;
aud[33264]=16'he4d3;
aud[33265]=16'he4e7;
aud[33266]=16'he4fa;
aud[33267]=16'he50e;
aud[33268]=16'he521;
aud[33269]=16'he535;
aud[33270]=16'he548;
aud[33271]=16'he55c;
aud[33272]=16'he56f;
aud[33273]=16'he583;
aud[33274]=16'he596;
aud[33275]=16'he5aa;
aud[33276]=16'he5bd;
aud[33277]=16'he5d1;
aud[33278]=16'he5e4;
aud[33279]=16'he5f8;
aud[33280]=16'he60c;
aud[33281]=16'he61f;
aud[33282]=16'he633;
aud[33283]=16'he646;
aud[33284]=16'he65a;
aud[33285]=16'he66e;
aud[33286]=16'he681;
aud[33287]=16'he695;
aud[33288]=16'he6a9;
aud[33289]=16'he6bd;
aud[33290]=16'he6d0;
aud[33291]=16'he6e4;
aud[33292]=16'he6f8;
aud[33293]=16'he70b;
aud[33294]=16'he71f;
aud[33295]=16'he733;
aud[33296]=16'he747;
aud[33297]=16'he75b;
aud[33298]=16'he76e;
aud[33299]=16'he782;
aud[33300]=16'he796;
aud[33301]=16'he7aa;
aud[33302]=16'he7be;
aud[33303]=16'he7d1;
aud[33304]=16'he7e5;
aud[33305]=16'he7f9;
aud[33306]=16'he80d;
aud[33307]=16'he821;
aud[33308]=16'he835;
aud[33309]=16'he849;
aud[33310]=16'he85d;
aud[33311]=16'he871;
aud[33312]=16'he885;
aud[33313]=16'he899;
aud[33314]=16'he8ad;
aud[33315]=16'he8c0;
aud[33316]=16'he8d4;
aud[33317]=16'he8e8;
aud[33318]=16'he8fc;
aud[33319]=16'he910;
aud[33320]=16'he925;
aud[33321]=16'he939;
aud[33322]=16'he94d;
aud[33323]=16'he961;
aud[33324]=16'he975;
aud[33325]=16'he989;
aud[33326]=16'he99d;
aud[33327]=16'he9b1;
aud[33328]=16'he9c5;
aud[33329]=16'he9d9;
aud[33330]=16'he9ed;
aud[33331]=16'hea01;
aud[33332]=16'hea16;
aud[33333]=16'hea2a;
aud[33334]=16'hea3e;
aud[33335]=16'hea52;
aud[33336]=16'hea66;
aud[33337]=16'hea7a;
aud[33338]=16'hea8f;
aud[33339]=16'heaa3;
aud[33340]=16'heab7;
aud[33341]=16'heacb;
aud[33342]=16'heae0;
aud[33343]=16'heaf4;
aud[33344]=16'heb08;
aud[33345]=16'heb1c;
aud[33346]=16'heb31;
aud[33347]=16'heb45;
aud[33348]=16'heb59;
aud[33349]=16'heb6e;
aud[33350]=16'heb82;
aud[33351]=16'heb96;
aud[33352]=16'hebab;
aud[33353]=16'hebbf;
aud[33354]=16'hebd3;
aud[33355]=16'hebe8;
aud[33356]=16'hebfc;
aud[33357]=16'hec10;
aud[33358]=16'hec25;
aud[33359]=16'hec39;
aud[33360]=16'hec4d;
aud[33361]=16'hec62;
aud[33362]=16'hec76;
aud[33363]=16'hec8b;
aud[33364]=16'hec9f;
aud[33365]=16'hecb4;
aud[33366]=16'hecc8;
aud[33367]=16'hecdd;
aud[33368]=16'hecf1;
aud[33369]=16'hed05;
aud[33370]=16'hed1a;
aud[33371]=16'hed2e;
aud[33372]=16'hed43;
aud[33373]=16'hed57;
aud[33374]=16'hed6c;
aud[33375]=16'hed81;
aud[33376]=16'hed95;
aud[33377]=16'hedaa;
aud[33378]=16'hedbe;
aud[33379]=16'hedd3;
aud[33380]=16'hede7;
aud[33381]=16'hedfc;
aud[33382]=16'hee10;
aud[33383]=16'hee25;
aud[33384]=16'hee3a;
aud[33385]=16'hee4e;
aud[33386]=16'hee63;
aud[33387]=16'hee77;
aud[33388]=16'hee8c;
aud[33389]=16'heea1;
aud[33390]=16'heeb5;
aud[33391]=16'heeca;
aud[33392]=16'heedf;
aud[33393]=16'heef3;
aud[33394]=16'hef08;
aud[33395]=16'hef1d;
aud[33396]=16'hef31;
aud[33397]=16'hef46;
aud[33398]=16'hef5b;
aud[33399]=16'hef70;
aud[33400]=16'hef84;
aud[33401]=16'hef99;
aud[33402]=16'hefae;
aud[33403]=16'hefc2;
aud[33404]=16'hefd7;
aud[33405]=16'hefec;
aud[33406]=16'hf001;
aud[33407]=16'hf015;
aud[33408]=16'hf02a;
aud[33409]=16'hf03f;
aud[33410]=16'hf054;
aud[33411]=16'hf069;
aud[33412]=16'hf07d;
aud[33413]=16'hf092;
aud[33414]=16'hf0a7;
aud[33415]=16'hf0bc;
aud[33416]=16'hf0d1;
aud[33417]=16'hf0e6;
aud[33418]=16'hf0fa;
aud[33419]=16'hf10f;
aud[33420]=16'hf124;
aud[33421]=16'hf139;
aud[33422]=16'hf14e;
aud[33423]=16'hf163;
aud[33424]=16'hf178;
aud[33425]=16'hf18c;
aud[33426]=16'hf1a1;
aud[33427]=16'hf1b6;
aud[33428]=16'hf1cb;
aud[33429]=16'hf1e0;
aud[33430]=16'hf1f5;
aud[33431]=16'hf20a;
aud[33432]=16'hf21f;
aud[33433]=16'hf234;
aud[33434]=16'hf249;
aud[33435]=16'hf25e;
aud[33436]=16'hf273;
aud[33437]=16'hf288;
aud[33438]=16'hf29d;
aud[33439]=16'hf2b2;
aud[33440]=16'hf2c7;
aud[33441]=16'hf2dc;
aud[33442]=16'hf2f1;
aud[33443]=16'hf306;
aud[33444]=16'hf31b;
aud[33445]=16'hf330;
aud[33446]=16'hf345;
aud[33447]=16'hf35a;
aud[33448]=16'hf36f;
aud[33449]=16'hf384;
aud[33450]=16'hf399;
aud[33451]=16'hf3ae;
aud[33452]=16'hf3c3;
aud[33453]=16'hf3d8;
aud[33454]=16'hf3ed;
aud[33455]=16'hf402;
aud[33456]=16'hf417;
aud[33457]=16'hf42c;
aud[33458]=16'hf441;
aud[33459]=16'hf456;
aud[33460]=16'hf46b;
aud[33461]=16'hf480;
aud[33462]=16'hf496;
aud[33463]=16'hf4ab;
aud[33464]=16'hf4c0;
aud[33465]=16'hf4d5;
aud[33466]=16'hf4ea;
aud[33467]=16'hf4ff;
aud[33468]=16'hf514;
aud[33469]=16'hf529;
aud[33470]=16'hf53f;
aud[33471]=16'hf554;
aud[33472]=16'hf569;
aud[33473]=16'hf57e;
aud[33474]=16'hf593;
aud[33475]=16'hf5a8;
aud[33476]=16'hf5bd;
aud[33477]=16'hf5d3;
aud[33478]=16'hf5e8;
aud[33479]=16'hf5fd;
aud[33480]=16'hf612;
aud[33481]=16'hf627;
aud[33482]=16'hf63d;
aud[33483]=16'hf652;
aud[33484]=16'hf667;
aud[33485]=16'hf67c;
aud[33486]=16'hf691;
aud[33487]=16'hf6a7;
aud[33488]=16'hf6bc;
aud[33489]=16'hf6d1;
aud[33490]=16'hf6e6;
aud[33491]=16'hf6fb;
aud[33492]=16'hf711;
aud[33493]=16'hf726;
aud[33494]=16'hf73b;
aud[33495]=16'hf750;
aud[33496]=16'hf766;
aud[33497]=16'hf77b;
aud[33498]=16'hf790;
aud[33499]=16'hf7a5;
aud[33500]=16'hf7bb;
aud[33501]=16'hf7d0;
aud[33502]=16'hf7e5;
aud[33503]=16'hf7fb;
aud[33504]=16'hf810;
aud[33505]=16'hf825;
aud[33506]=16'hf83a;
aud[33507]=16'hf850;
aud[33508]=16'hf865;
aud[33509]=16'hf87a;
aud[33510]=16'hf890;
aud[33511]=16'hf8a5;
aud[33512]=16'hf8ba;
aud[33513]=16'hf8cf;
aud[33514]=16'hf8e5;
aud[33515]=16'hf8fa;
aud[33516]=16'hf90f;
aud[33517]=16'hf925;
aud[33518]=16'hf93a;
aud[33519]=16'hf94f;
aud[33520]=16'hf965;
aud[33521]=16'hf97a;
aud[33522]=16'hf98f;
aud[33523]=16'hf9a5;
aud[33524]=16'hf9ba;
aud[33525]=16'hf9cf;
aud[33526]=16'hf9e5;
aud[33527]=16'hf9fa;
aud[33528]=16'hfa0f;
aud[33529]=16'hfa25;
aud[33530]=16'hfa3a;
aud[33531]=16'hfa50;
aud[33532]=16'hfa65;
aud[33533]=16'hfa7a;
aud[33534]=16'hfa90;
aud[33535]=16'hfaa5;
aud[33536]=16'hfaba;
aud[33537]=16'hfad0;
aud[33538]=16'hfae5;
aud[33539]=16'hfafb;
aud[33540]=16'hfb10;
aud[33541]=16'hfb25;
aud[33542]=16'hfb3b;
aud[33543]=16'hfb50;
aud[33544]=16'hfb65;
aud[33545]=16'hfb7b;
aud[33546]=16'hfb90;
aud[33547]=16'hfba6;
aud[33548]=16'hfbbb;
aud[33549]=16'hfbd0;
aud[33550]=16'hfbe6;
aud[33551]=16'hfbfb;
aud[33552]=16'hfc11;
aud[33553]=16'hfc26;
aud[33554]=16'hfc3b;
aud[33555]=16'hfc51;
aud[33556]=16'hfc66;
aud[33557]=16'hfc7c;
aud[33558]=16'hfc91;
aud[33559]=16'hfca7;
aud[33560]=16'hfcbc;
aud[33561]=16'hfcd1;
aud[33562]=16'hfce7;
aud[33563]=16'hfcfc;
aud[33564]=16'hfd12;
aud[33565]=16'hfd27;
aud[33566]=16'hfd3c;
aud[33567]=16'hfd52;
aud[33568]=16'hfd67;
aud[33569]=16'hfd7d;
aud[33570]=16'hfd92;
aud[33571]=16'hfda8;
aud[33572]=16'hfdbd;
aud[33573]=16'hfdd2;
aud[33574]=16'hfde8;
aud[33575]=16'hfdfd;
aud[33576]=16'hfe13;
aud[33577]=16'hfe28;
aud[33578]=16'hfe3e;
aud[33579]=16'hfe53;
aud[33580]=16'hfe69;
aud[33581]=16'hfe7e;
aud[33582]=16'hfe93;
aud[33583]=16'hfea9;
aud[33584]=16'hfebe;
aud[33585]=16'hfed4;
aud[33586]=16'hfee9;
aud[33587]=16'hfeff;
aud[33588]=16'hff14;
aud[33589]=16'hff2a;
aud[33590]=16'hff3f;
aud[33591]=16'hff54;
aud[33592]=16'hff6a;
aud[33593]=16'hff7f;
aud[33594]=16'hff95;
aud[33595]=16'hffaa;
aud[33596]=16'hffc0;
aud[33597]=16'hffd5;
aud[33598]=16'hffeb;
aud[33599]=16'h0;
aud[33600]=16'h15;
aud[33601]=16'h2b;
aud[33602]=16'h40;
aud[33603]=16'h56;
aud[33604]=16'h6b;
aud[33605]=16'h81;
aud[33606]=16'h96;
aud[33607]=16'hac;
aud[33608]=16'hc1;
aud[33609]=16'hd6;
aud[33610]=16'hec;
aud[33611]=16'h101;
aud[33612]=16'h117;
aud[33613]=16'h12c;
aud[33614]=16'h142;
aud[33615]=16'h157;
aud[33616]=16'h16d;
aud[33617]=16'h182;
aud[33618]=16'h197;
aud[33619]=16'h1ad;
aud[33620]=16'h1c2;
aud[33621]=16'h1d8;
aud[33622]=16'h1ed;
aud[33623]=16'h203;
aud[33624]=16'h218;
aud[33625]=16'h22e;
aud[33626]=16'h243;
aud[33627]=16'h258;
aud[33628]=16'h26e;
aud[33629]=16'h283;
aud[33630]=16'h299;
aud[33631]=16'h2ae;
aud[33632]=16'h2c4;
aud[33633]=16'h2d9;
aud[33634]=16'h2ee;
aud[33635]=16'h304;
aud[33636]=16'h319;
aud[33637]=16'h32f;
aud[33638]=16'h344;
aud[33639]=16'h359;
aud[33640]=16'h36f;
aud[33641]=16'h384;
aud[33642]=16'h39a;
aud[33643]=16'h3af;
aud[33644]=16'h3c5;
aud[33645]=16'h3da;
aud[33646]=16'h3ef;
aud[33647]=16'h405;
aud[33648]=16'h41a;
aud[33649]=16'h430;
aud[33650]=16'h445;
aud[33651]=16'h45a;
aud[33652]=16'h470;
aud[33653]=16'h485;
aud[33654]=16'h49b;
aud[33655]=16'h4b0;
aud[33656]=16'h4c5;
aud[33657]=16'h4db;
aud[33658]=16'h4f0;
aud[33659]=16'h505;
aud[33660]=16'h51b;
aud[33661]=16'h530;
aud[33662]=16'h546;
aud[33663]=16'h55b;
aud[33664]=16'h570;
aud[33665]=16'h586;
aud[33666]=16'h59b;
aud[33667]=16'h5b0;
aud[33668]=16'h5c6;
aud[33669]=16'h5db;
aud[33670]=16'h5f1;
aud[33671]=16'h606;
aud[33672]=16'h61b;
aud[33673]=16'h631;
aud[33674]=16'h646;
aud[33675]=16'h65b;
aud[33676]=16'h671;
aud[33677]=16'h686;
aud[33678]=16'h69b;
aud[33679]=16'h6b1;
aud[33680]=16'h6c6;
aud[33681]=16'h6db;
aud[33682]=16'h6f1;
aud[33683]=16'h706;
aud[33684]=16'h71b;
aud[33685]=16'h731;
aud[33686]=16'h746;
aud[33687]=16'h75b;
aud[33688]=16'h770;
aud[33689]=16'h786;
aud[33690]=16'h79b;
aud[33691]=16'h7b0;
aud[33692]=16'h7c6;
aud[33693]=16'h7db;
aud[33694]=16'h7f0;
aud[33695]=16'h805;
aud[33696]=16'h81b;
aud[33697]=16'h830;
aud[33698]=16'h845;
aud[33699]=16'h85b;
aud[33700]=16'h870;
aud[33701]=16'h885;
aud[33702]=16'h89a;
aud[33703]=16'h8b0;
aud[33704]=16'h8c5;
aud[33705]=16'h8da;
aud[33706]=16'h8ef;
aud[33707]=16'h905;
aud[33708]=16'h91a;
aud[33709]=16'h92f;
aud[33710]=16'h944;
aud[33711]=16'h959;
aud[33712]=16'h96f;
aud[33713]=16'h984;
aud[33714]=16'h999;
aud[33715]=16'h9ae;
aud[33716]=16'h9c3;
aud[33717]=16'h9d9;
aud[33718]=16'h9ee;
aud[33719]=16'ha03;
aud[33720]=16'ha18;
aud[33721]=16'ha2d;
aud[33722]=16'ha43;
aud[33723]=16'ha58;
aud[33724]=16'ha6d;
aud[33725]=16'ha82;
aud[33726]=16'ha97;
aud[33727]=16'haac;
aud[33728]=16'hac1;
aud[33729]=16'had7;
aud[33730]=16'haec;
aud[33731]=16'hb01;
aud[33732]=16'hb16;
aud[33733]=16'hb2b;
aud[33734]=16'hb40;
aud[33735]=16'hb55;
aud[33736]=16'hb6a;
aud[33737]=16'hb80;
aud[33738]=16'hb95;
aud[33739]=16'hbaa;
aud[33740]=16'hbbf;
aud[33741]=16'hbd4;
aud[33742]=16'hbe9;
aud[33743]=16'hbfe;
aud[33744]=16'hc13;
aud[33745]=16'hc28;
aud[33746]=16'hc3d;
aud[33747]=16'hc52;
aud[33748]=16'hc67;
aud[33749]=16'hc7c;
aud[33750]=16'hc91;
aud[33751]=16'hca6;
aud[33752]=16'hcbb;
aud[33753]=16'hcd0;
aud[33754]=16'hce5;
aud[33755]=16'hcfa;
aud[33756]=16'hd0f;
aud[33757]=16'hd24;
aud[33758]=16'hd39;
aud[33759]=16'hd4e;
aud[33760]=16'hd63;
aud[33761]=16'hd78;
aud[33762]=16'hd8d;
aud[33763]=16'hda2;
aud[33764]=16'hdb7;
aud[33765]=16'hdcc;
aud[33766]=16'hde1;
aud[33767]=16'hdf6;
aud[33768]=16'he0b;
aud[33769]=16'he20;
aud[33770]=16'he35;
aud[33771]=16'he4a;
aud[33772]=16'he5f;
aud[33773]=16'he74;
aud[33774]=16'he88;
aud[33775]=16'he9d;
aud[33776]=16'heb2;
aud[33777]=16'hec7;
aud[33778]=16'hedc;
aud[33779]=16'hef1;
aud[33780]=16'hf06;
aud[33781]=16'hf1a;
aud[33782]=16'hf2f;
aud[33783]=16'hf44;
aud[33784]=16'hf59;
aud[33785]=16'hf6e;
aud[33786]=16'hf83;
aud[33787]=16'hf97;
aud[33788]=16'hfac;
aud[33789]=16'hfc1;
aud[33790]=16'hfd6;
aud[33791]=16'hfeb;
aud[33792]=16'hfff;
aud[33793]=16'h1014;
aud[33794]=16'h1029;
aud[33795]=16'h103e;
aud[33796]=16'h1052;
aud[33797]=16'h1067;
aud[33798]=16'h107c;
aud[33799]=16'h1090;
aud[33800]=16'h10a5;
aud[33801]=16'h10ba;
aud[33802]=16'h10cf;
aud[33803]=16'h10e3;
aud[33804]=16'h10f8;
aud[33805]=16'h110d;
aud[33806]=16'h1121;
aud[33807]=16'h1136;
aud[33808]=16'h114b;
aud[33809]=16'h115f;
aud[33810]=16'h1174;
aud[33811]=16'h1189;
aud[33812]=16'h119d;
aud[33813]=16'h11b2;
aud[33814]=16'h11c6;
aud[33815]=16'h11db;
aud[33816]=16'h11f0;
aud[33817]=16'h1204;
aud[33818]=16'h1219;
aud[33819]=16'h122d;
aud[33820]=16'h1242;
aud[33821]=16'h1256;
aud[33822]=16'h126b;
aud[33823]=16'h127f;
aud[33824]=16'h1294;
aud[33825]=16'h12a9;
aud[33826]=16'h12bd;
aud[33827]=16'h12d2;
aud[33828]=16'h12e6;
aud[33829]=16'h12fb;
aud[33830]=16'h130f;
aud[33831]=16'h1323;
aud[33832]=16'h1338;
aud[33833]=16'h134c;
aud[33834]=16'h1361;
aud[33835]=16'h1375;
aud[33836]=16'h138a;
aud[33837]=16'h139e;
aud[33838]=16'h13b3;
aud[33839]=16'h13c7;
aud[33840]=16'h13db;
aud[33841]=16'h13f0;
aud[33842]=16'h1404;
aud[33843]=16'h1418;
aud[33844]=16'h142d;
aud[33845]=16'h1441;
aud[33846]=16'h1455;
aud[33847]=16'h146a;
aud[33848]=16'h147e;
aud[33849]=16'h1492;
aud[33850]=16'h14a7;
aud[33851]=16'h14bb;
aud[33852]=16'h14cf;
aud[33853]=16'h14e4;
aud[33854]=16'h14f8;
aud[33855]=16'h150c;
aud[33856]=16'h1520;
aud[33857]=16'h1535;
aud[33858]=16'h1549;
aud[33859]=16'h155d;
aud[33860]=16'h1571;
aud[33861]=16'h1586;
aud[33862]=16'h159a;
aud[33863]=16'h15ae;
aud[33864]=16'h15c2;
aud[33865]=16'h15d6;
aud[33866]=16'h15ea;
aud[33867]=16'h15ff;
aud[33868]=16'h1613;
aud[33869]=16'h1627;
aud[33870]=16'h163b;
aud[33871]=16'h164f;
aud[33872]=16'h1663;
aud[33873]=16'h1677;
aud[33874]=16'h168b;
aud[33875]=16'h169f;
aud[33876]=16'h16b3;
aud[33877]=16'h16c7;
aud[33878]=16'h16db;
aud[33879]=16'h16f0;
aud[33880]=16'h1704;
aud[33881]=16'h1718;
aud[33882]=16'h172c;
aud[33883]=16'h1740;
aud[33884]=16'h1753;
aud[33885]=16'h1767;
aud[33886]=16'h177b;
aud[33887]=16'h178f;
aud[33888]=16'h17a3;
aud[33889]=16'h17b7;
aud[33890]=16'h17cb;
aud[33891]=16'h17df;
aud[33892]=16'h17f3;
aud[33893]=16'h1807;
aud[33894]=16'h181b;
aud[33895]=16'h182f;
aud[33896]=16'h1842;
aud[33897]=16'h1856;
aud[33898]=16'h186a;
aud[33899]=16'h187e;
aud[33900]=16'h1892;
aud[33901]=16'h18a5;
aud[33902]=16'h18b9;
aud[33903]=16'h18cd;
aud[33904]=16'h18e1;
aud[33905]=16'h18f5;
aud[33906]=16'h1908;
aud[33907]=16'h191c;
aud[33908]=16'h1930;
aud[33909]=16'h1943;
aud[33910]=16'h1957;
aud[33911]=16'h196b;
aud[33912]=16'h197f;
aud[33913]=16'h1992;
aud[33914]=16'h19a6;
aud[33915]=16'h19ba;
aud[33916]=16'h19cd;
aud[33917]=16'h19e1;
aud[33918]=16'h19f4;
aud[33919]=16'h1a08;
aud[33920]=16'h1a1c;
aud[33921]=16'h1a2f;
aud[33922]=16'h1a43;
aud[33923]=16'h1a56;
aud[33924]=16'h1a6a;
aud[33925]=16'h1a7d;
aud[33926]=16'h1a91;
aud[33927]=16'h1aa4;
aud[33928]=16'h1ab8;
aud[33929]=16'h1acb;
aud[33930]=16'h1adf;
aud[33931]=16'h1af2;
aud[33932]=16'h1b06;
aud[33933]=16'h1b19;
aud[33934]=16'h1b2d;
aud[33935]=16'h1b40;
aud[33936]=16'h1b53;
aud[33937]=16'h1b67;
aud[33938]=16'h1b7a;
aud[33939]=16'h1b8d;
aud[33940]=16'h1ba1;
aud[33941]=16'h1bb4;
aud[33942]=16'h1bc8;
aud[33943]=16'h1bdb;
aud[33944]=16'h1bee;
aud[33945]=16'h1c01;
aud[33946]=16'h1c15;
aud[33947]=16'h1c28;
aud[33948]=16'h1c3b;
aud[33949]=16'h1c4e;
aud[33950]=16'h1c62;
aud[33951]=16'h1c75;
aud[33952]=16'h1c88;
aud[33953]=16'h1c9b;
aud[33954]=16'h1cae;
aud[33955]=16'h1cc2;
aud[33956]=16'h1cd5;
aud[33957]=16'h1ce8;
aud[33958]=16'h1cfb;
aud[33959]=16'h1d0e;
aud[33960]=16'h1d21;
aud[33961]=16'h1d34;
aud[33962]=16'h1d47;
aud[33963]=16'h1d5b;
aud[33964]=16'h1d6e;
aud[33965]=16'h1d81;
aud[33966]=16'h1d94;
aud[33967]=16'h1da7;
aud[33968]=16'h1dba;
aud[33969]=16'h1dcd;
aud[33970]=16'h1de0;
aud[33971]=16'h1df3;
aud[33972]=16'h1e06;
aud[33973]=16'h1e18;
aud[33974]=16'h1e2b;
aud[33975]=16'h1e3e;
aud[33976]=16'h1e51;
aud[33977]=16'h1e64;
aud[33978]=16'h1e77;
aud[33979]=16'h1e8a;
aud[33980]=16'h1e9d;
aud[33981]=16'h1eaf;
aud[33982]=16'h1ec2;
aud[33983]=16'h1ed5;
aud[33984]=16'h1ee8;
aud[33985]=16'h1efb;
aud[33986]=16'h1f0d;
aud[33987]=16'h1f20;
aud[33988]=16'h1f33;
aud[33989]=16'h1f46;
aud[33990]=16'h1f58;
aud[33991]=16'h1f6b;
aud[33992]=16'h1f7e;
aud[33993]=16'h1f90;
aud[33994]=16'h1fa3;
aud[33995]=16'h1fb6;
aud[33996]=16'h1fc8;
aud[33997]=16'h1fdb;
aud[33998]=16'h1fed;
aud[33999]=16'h2000;
aud[34000]=16'h2013;
aud[34001]=16'h2025;
aud[34002]=16'h2038;
aud[34003]=16'h204a;
aud[34004]=16'h205d;
aud[34005]=16'h206f;
aud[34006]=16'h2082;
aud[34007]=16'h2094;
aud[34008]=16'h20a7;
aud[34009]=16'h20b9;
aud[34010]=16'h20cb;
aud[34011]=16'h20de;
aud[34012]=16'h20f0;
aud[34013]=16'h2103;
aud[34014]=16'h2115;
aud[34015]=16'h2127;
aud[34016]=16'h213a;
aud[34017]=16'h214c;
aud[34018]=16'h215e;
aud[34019]=16'h2171;
aud[34020]=16'h2183;
aud[34021]=16'h2195;
aud[34022]=16'h21a7;
aud[34023]=16'h21ba;
aud[34024]=16'h21cc;
aud[34025]=16'h21de;
aud[34026]=16'h21f0;
aud[34027]=16'h2202;
aud[34028]=16'h2215;
aud[34029]=16'h2227;
aud[34030]=16'h2239;
aud[34031]=16'h224b;
aud[34032]=16'h225d;
aud[34033]=16'h226f;
aud[34034]=16'h2281;
aud[34035]=16'h2293;
aud[34036]=16'h22a5;
aud[34037]=16'h22b7;
aud[34038]=16'h22c9;
aud[34039]=16'h22db;
aud[34040]=16'h22ed;
aud[34041]=16'h22ff;
aud[34042]=16'h2311;
aud[34043]=16'h2323;
aud[34044]=16'h2335;
aud[34045]=16'h2347;
aud[34046]=16'h2359;
aud[34047]=16'h236b;
aud[34048]=16'h237d;
aud[34049]=16'h238e;
aud[34050]=16'h23a0;
aud[34051]=16'h23b2;
aud[34052]=16'h23c4;
aud[34053]=16'h23d6;
aud[34054]=16'h23e7;
aud[34055]=16'h23f9;
aud[34056]=16'h240b;
aud[34057]=16'h241d;
aud[34058]=16'h242e;
aud[34059]=16'h2440;
aud[34060]=16'h2452;
aud[34061]=16'h2463;
aud[34062]=16'h2475;
aud[34063]=16'h2487;
aud[34064]=16'h2498;
aud[34065]=16'h24aa;
aud[34066]=16'h24bb;
aud[34067]=16'h24cd;
aud[34068]=16'h24de;
aud[34069]=16'h24f0;
aud[34070]=16'h2501;
aud[34071]=16'h2513;
aud[34072]=16'h2524;
aud[34073]=16'h2536;
aud[34074]=16'h2547;
aud[34075]=16'h2559;
aud[34076]=16'h256a;
aud[34077]=16'h257c;
aud[34078]=16'h258d;
aud[34079]=16'h259e;
aud[34080]=16'h25b0;
aud[34081]=16'h25c1;
aud[34082]=16'h25d2;
aud[34083]=16'h25e4;
aud[34084]=16'h25f5;
aud[34085]=16'h2606;
aud[34086]=16'h2617;
aud[34087]=16'h2629;
aud[34088]=16'h263a;
aud[34089]=16'h264b;
aud[34090]=16'h265c;
aud[34091]=16'h266d;
aud[34092]=16'h267e;
aud[34093]=16'h2690;
aud[34094]=16'h26a1;
aud[34095]=16'h26b2;
aud[34096]=16'h26c3;
aud[34097]=16'h26d4;
aud[34098]=16'h26e5;
aud[34099]=16'h26f6;
aud[34100]=16'h2707;
aud[34101]=16'h2718;
aud[34102]=16'h2729;
aud[34103]=16'h273a;
aud[34104]=16'h274b;
aud[34105]=16'h275c;
aud[34106]=16'h276d;
aud[34107]=16'h277e;
aud[34108]=16'h278e;
aud[34109]=16'h279f;
aud[34110]=16'h27b0;
aud[34111]=16'h27c1;
aud[34112]=16'h27d2;
aud[34113]=16'h27e2;
aud[34114]=16'h27f3;
aud[34115]=16'h2804;
aud[34116]=16'h2815;
aud[34117]=16'h2825;
aud[34118]=16'h2836;
aud[34119]=16'h2847;
aud[34120]=16'h2857;
aud[34121]=16'h2868;
aud[34122]=16'h2879;
aud[34123]=16'h2889;
aud[34124]=16'h289a;
aud[34125]=16'h28aa;
aud[34126]=16'h28bb;
aud[34127]=16'h28cc;
aud[34128]=16'h28dc;
aud[34129]=16'h28ed;
aud[34130]=16'h28fd;
aud[34131]=16'h290e;
aud[34132]=16'h291e;
aud[34133]=16'h292e;
aud[34134]=16'h293f;
aud[34135]=16'h294f;
aud[34136]=16'h2960;
aud[34137]=16'h2970;
aud[34138]=16'h2980;
aud[34139]=16'h2991;
aud[34140]=16'h29a1;
aud[34141]=16'h29b1;
aud[34142]=16'h29c1;
aud[34143]=16'h29d2;
aud[34144]=16'h29e2;
aud[34145]=16'h29f2;
aud[34146]=16'h2a02;
aud[34147]=16'h2a12;
aud[34148]=16'h2a23;
aud[34149]=16'h2a33;
aud[34150]=16'h2a43;
aud[34151]=16'h2a53;
aud[34152]=16'h2a63;
aud[34153]=16'h2a73;
aud[34154]=16'h2a83;
aud[34155]=16'h2a93;
aud[34156]=16'h2aa3;
aud[34157]=16'h2ab3;
aud[34158]=16'h2ac3;
aud[34159]=16'h2ad3;
aud[34160]=16'h2ae3;
aud[34161]=16'h2af3;
aud[34162]=16'h2b03;
aud[34163]=16'h2b13;
aud[34164]=16'h2b22;
aud[34165]=16'h2b32;
aud[34166]=16'h2b42;
aud[34167]=16'h2b52;
aud[34168]=16'h2b62;
aud[34169]=16'h2b71;
aud[34170]=16'h2b81;
aud[34171]=16'h2b91;
aud[34172]=16'h2ba1;
aud[34173]=16'h2bb0;
aud[34174]=16'h2bc0;
aud[34175]=16'h2bd0;
aud[34176]=16'h2bdf;
aud[34177]=16'h2bef;
aud[34178]=16'h2bfe;
aud[34179]=16'h2c0e;
aud[34180]=16'h2c1e;
aud[34181]=16'h2c2d;
aud[34182]=16'h2c3d;
aud[34183]=16'h2c4c;
aud[34184]=16'h2c5c;
aud[34185]=16'h2c6b;
aud[34186]=16'h2c7a;
aud[34187]=16'h2c8a;
aud[34188]=16'h2c99;
aud[34189]=16'h2ca9;
aud[34190]=16'h2cb8;
aud[34191]=16'h2cc7;
aud[34192]=16'h2cd7;
aud[34193]=16'h2ce6;
aud[34194]=16'h2cf5;
aud[34195]=16'h2d04;
aud[34196]=16'h2d14;
aud[34197]=16'h2d23;
aud[34198]=16'h2d32;
aud[34199]=16'h2d41;
aud[34200]=16'h2d50;
aud[34201]=16'h2d60;
aud[34202]=16'h2d6f;
aud[34203]=16'h2d7e;
aud[34204]=16'h2d8d;
aud[34205]=16'h2d9c;
aud[34206]=16'h2dab;
aud[34207]=16'h2dba;
aud[34208]=16'h2dc9;
aud[34209]=16'h2dd8;
aud[34210]=16'h2de7;
aud[34211]=16'h2df6;
aud[34212]=16'h2e05;
aud[34213]=16'h2e14;
aud[34214]=16'h2e22;
aud[34215]=16'h2e31;
aud[34216]=16'h2e40;
aud[34217]=16'h2e4f;
aud[34218]=16'h2e5e;
aud[34219]=16'h2e6d;
aud[34220]=16'h2e7b;
aud[34221]=16'h2e8a;
aud[34222]=16'h2e99;
aud[34223]=16'h2ea7;
aud[34224]=16'h2eb6;
aud[34225]=16'h2ec5;
aud[34226]=16'h2ed3;
aud[34227]=16'h2ee2;
aud[34228]=16'h2ef1;
aud[34229]=16'h2eff;
aud[34230]=16'h2f0e;
aud[34231]=16'h2f1c;
aud[34232]=16'h2f2b;
aud[34233]=16'h2f39;
aud[34234]=16'h2f48;
aud[34235]=16'h2f56;
aud[34236]=16'h2f65;
aud[34237]=16'h2f73;
aud[34238]=16'h2f81;
aud[34239]=16'h2f90;
aud[34240]=16'h2f9e;
aud[34241]=16'h2fac;
aud[34242]=16'h2fbb;
aud[34243]=16'h2fc9;
aud[34244]=16'h2fd7;
aud[34245]=16'h2fe5;
aud[34246]=16'h2ff4;
aud[34247]=16'h3002;
aud[34248]=16'h3010;
aud[34249]=16'h301e;
aud[34250]=16'h302c;
aud[34251]=16'h303a;
aud[34252]=16'h3048;
aud[34253]=16'h3057;
aud[34254]=16'h3065;
aud[34255]=16'h3073;
aud[34256]=16'h3081;
aud[34257]=16'h308f;
aud[34258]=16'h309d;
aud[34259]=16'h30aa;
aud[34260]=16'h30b8;
aud[34261]=16'h30c6;
aud[34262]=16'h30d4;
aud[34263]=16'h30e2;
aud[34264]=16'h30f0;
aud[34265]=16'h30fe;
aud[34266]=16'h310b;
aud[34267]=16'h3119;
aud[34268]=16'h3127;
aud[34269]=16'h3135;
aud[34270]=16'h3142;
aud[34271]=16'h3150;
aud[34272]=16'h315e;
aud[34273]=16'h316b;
aud[34274]=16'h3179;
aud[34275]=16'h3187;
aud[34276]=16'h3194;
aud[34277]=16'h31a2;
aud[34278]=16'h31af;
aud[34279]=16'h31bd;
aud[34280]=16'h31ca;
aud[34281]=16'h31d8;
aud[34282]=16'h31e5;
aud[34283]=16'h31f3;
aud[34284]=16'h3200;
aud[34285]=16'h320d;
aud[34286]=16'h321b;
aud[34287]=16'h3228;
aud[34288]=16'h3235;
aud[34289]=16'h3243;
aud[34290]=16'h3250;
aud[34291]=16'h325d;
aud[34292]=16'h326a;
aud[34293]=16'h3278;
aud[34294]=16'h3285;
aud[34295]=16'h3292;
aud[34296]=16'h329f;
aud[34297]=16'h32ac;
aud[34298]=16'h32b9;
aud[34299]=16'h32c6;
aud[34300]=16'h32d3;
aud[34301]=16'h32e0;
aud[34302]=16'h32ed;
aud[34303]=16'h32fa;
aud[34304]=16'h3307;
aud[34305]=16'h3314;
aud[34306]=16'h3321;
aud[34307]=16'h332e;
aud[34308]=16'h333b;
aud[34309]=16'h3348;
aud[34310]=16'h3355;
aud[34311]=16'h3361;
aud[34312]=16'h336e;
aud[34313]=16'h337b;
aud[34314]=16'h3388;
aud[34315]=16'h3394;
aud[34316]=16'h33a1;
aud[34317]=16'h33ae;
aud[34318]=16'h33ba;
aud[34319]=16'h33c7;
aud[34320]=16'h33d4;
aud[34321]=16'h33e0;
aud[34322]=16'h33ed;
aud[34323]=16'h33f9;
aud[34324]=16'h3406;
aud[34325]=16'h3412;
aud[34326]=16'h341f;
aud[34327]=16'h342b;
aud[34328]=16'h3437;
aud[34329]=16'h3444;
aud[34330]=16'h3450;
aud[34331]=16'h345d;
aud[34332]=16'h3469;
aud[34333]=16'h3475;
aud[34334]=16'h3481;
aud[34335]=16'h348e;
aud[34336]=16'h349a;
aud[34337]=16'h34a6;
aud[34338]=16'h34b2;
aud[34339]=16'h34be;
aud[34340]=16'h34cb;
aud[34341]=16'h34d7;
aud[34342]=16'h34e3;
aud[34343]=16'h34ef;
aud[34344]=16'h34fb;
aud[34345]=16'h3507;
aud[34346]=16'h3513;
aud[34347]=16'h351f;
aud[34348]=16'h352b;
aud[34349]=16'h3537;
aud[34350]=16'h3543;
aud[34351]=16'h354f;
aud[34352]=16'h355a;
aud[34353]=16'h3566;
aud[34354]=16'h3572;
aud[34355]=16'h357e;
aud[34356]=16'h358a;
aud[34357]=16'h3595;
aud[34358]=16'h35a1;
aud[34359]=16'h35ad;
aud[34360]=16'h35b8;
aud[34361]=16'h35c4;
aud[34362]=16'h35d0;
aud[34363]=16'h35db;
aud[34364]=16'h35e7;
aud[34365]=16'h35f2;
aud[34366]=16'h35fe;
aud[34367]=16'h3609;
aud[34368]=16'h3615;
aud[34369]=16'h3620;
aud[34370]=16'h362c;
aud[34371]=16'h3637;
aud[34372]=16'h3643;
aud[34373]=16'h364e;
aud[34374]=16'h3659;
aud[34375]=16'h3665;
aud[34376]=16'h3670;
aud[34377]=16'h367b;
aud[34378]=16'h3686;
aud[34379]=16'h3692;
aud[34380]=16'h369d;
aud[34381]=16'h36a8;
aud[34382]=16'h36b3;
aud[34383]=16'h36be;
aud[34384]=16'h36c9;
aud[34385]=16'h36d4;
aud[34386]=16'h36e0;
aud[34387]=16'h36eb;
aud[34388]=16'h36f6;
aud[34389]=16'h3701;
aud[34390]=16'h370b;
aud[34391]=16'h3716;
aud[34392]=16'h3721;
aud[34393]=16'h372c;
aud[34394]=16'h3737;
aud[34395]=16'h3742;
aud[34396]=16'h374d;
aud[34397]=16'h3757;
aud[34398]=16'h3762;
aud[34399]=16'h376d;
aud[34400]=16'h3778;
aud[34401]=16'h3782;
aud[34402]=16'h378d;
aud[34403]=16'h3798;
aud[34404]=16'h37a2;
aud[34405]=16'h37ad;
aud[34406]=16'h37b7;
aud[34407]=16'h37c2;
aud[34408]=16'h37cc;
aud[34409]=16'h37d7;
aud[34410]=16'h37e1;
aud[34411]=16'h37ec;
aud[34412]=16'h37f6;
aud[34413]=16'h3801;
aud[34414]=16'h380b;
aud[34415]=16'h3815;
aud[34416]=16'h3820;
aud[34417]=16'h382a;
aud[34418]=16'h3834;
aud[34419]=16'h383f;
aud[34420]=16'h3849;
aud[34421]=16'h3853;
aud[34422]=16'h385d;
aud[34423]=16'h3867;
aud[34424]=16'h3871;
aud[34425]=16'h387b;
aud[34426]=16'h3886;
aud[34427]=16'h3890;
aud[34428]=16'h389a;
aud[34429]=16'h38a4;
aud[34430]=16'h38ae;
aud[34431]=16'h38b8;
aud[34432]=16'h38c1;
aud[34433]=16'h38cb;
aud[34434]=16'h38d5;
aud[34435]=16'h38df;
aud[34436]=16'h38e9;
aud[34437]=16'h38f3;
aud[34438]=16'h38fd;
aud[34439]=16'h3906;
aud[34440]=16'h3910;
aud[34441]=16'h391a;
aud[34442]=16'h3923;
aud[34443]=16'h392d;
aud[34444]=16'h3937;
aud[34445]=16'h3940;
aud[34446]=16'h394a;
aud[34447]=16'h3953;
aud[34448]=16'h395d;
aud[34449]=16'h3966;
aud[34450]=16'h3970;
aud[34451]=16'h3979;
aud[34452]=16'h3983;
aud[34453]=16'h398c;
aud[34454]=16'h3995;
aud[34455]=16'h399f;
aud[34456]=16'h39a8;
aud[34457]=16'h39b1;
aud[34458]=16'h39bb;
aud[34459]=16'h39c4;
aud[34460]=16'h39cd;
aud[34461]=16'h39d6;
aud[34462]=16'h39e0;
aud[34463]=16'h39e9;
aud[34464]=16'h39f2;
aud[34465]=16'h39fb;
aud[34466]=16'h3a04;
aud[34467]=16'h3a0d;
aud[34468]=16'h3a16;
aud[34469]=16'h3a1f;
aud[34470]=16'h3a28;
aud[34471]=16'h3a31;
aud[34472]=16'h3a3a;
aud[34473]=16'h3a43;
aud[34474]=16'h3a4c;
aud[34475]=16'h3a54;
aud[34476]=16'h3a5d;
aud[34477]=16'h3a66;
aud[34478]=16'h3a6f;
aud[34479]=16'h3a78;
aud[34480]=16'h3a80;
aud[34481]=16'h3a89;
aud[34482]=16'h3a92;
aud[34483]=16'h3a9a;
aud[34484]=16'h3aa3;
aud[34485]=16'h3aab;
aud[34486]=16'h3ab4;
aud[34487]=16'h3abc;
aud[34488]=16'h3ac5;
aud[34489]=16'h3acd;
aud[34490]=16'h3ad6;
aud[34491]=16'h3ade;
aud[34492]=16'h3ae7;
aud[34493]=16'h3aef;
aud[34494]=16'h3af7;
aud[34495]=16'h3b00;
aud[34496]=16'h3b08;
aud[34497]=16'h3b10;
aud[34498]=16'h3b19;
aud[34499]=16'h3b21;
aud[34500]=16'h3b29;
aud[34501]=16'h3b31;
aud[34502]=16'h3b39;
aud[34503]=16'h3b41;
aud[34504]=16'h3b4a;
aud[34505]=16'h3b52;
aud[34506]=16'h3b5a;
aud[34507]=16'h3b62;
aud[34508]=16'h3b6a;
aud[34509]=16'h3b72;
aud[34510]=16'h3b7a;
aud[34511]=16'h3b81;
aud[34512]=16'h3b89;
aud[34513]=16'h3b91;
aud[34514]=16'h3b99;
aud[34515]=16'h3ba1;
aud[34516]=16'h3ba9;
aud[34517]=16'h3bb0;
aud[34518]=16'h3bb8;
aud[34519]=16'h3bc0;
aud[34520]=16'h3bc7;
aud[34521]=16'h3bcf;
aud[34522]=16'h3bd7;
aud[34523]=16'h3bde;
aud[34524]=16'h3be6;
aud[34525]=16'h3bed;
aud[34526]=16'h3bf5;
aud[34527]=16'h3bfc;
aud[34528]=16'h3c04;
aud[34529]=16'h3c0b;
aud[34530]=16'h3c13;
aud[34531]=16'h3c1a;
aud[34532]=16'h3c21;
aud[34533]=16'h3c29;
aud[34534]=16'h3c30;
aud[34535]=16'h3c37;
aud[34536]=16'h3c3f;
aud[34537]=16'h3c46;
aud[34538]=16'h3c4d;
aud[34539]=16'h3c54;
aud[34540]=16'h3c5b;
aud[34541]=16'h3c63;
aud[34542]=16'h3c6a;
aud[34543]=16'h3c71;
aud[34544]=16'h3c78;
aud[34545]=16'h3c7f;
aud[34546]=16'h3c86;
aud[34547]=16'h3c8d;
aud[34548]=16'h3c94;
aud[34549]=16'h3c9b;
aud[34550]=16'h3ca1;
aud[34551]=16'h3ca8;
aud[34552]=16'h3caf;
aud[34553]=16'h3cb6;
aud[34554]=16'h3cbd;
aud[34555]=16'h3cc3;
aud[34556]=16'h3cca;
aud[34557]=16'h3cd1;
aud[34558]=16'h3cd7;
aud[34559]=16'h3cde;
aud[34560]=16'h3ce5;
aud[34561]=16'h3ceb;
aud[34562]=16'h3cf2;
aud[34563]=16'h3cf8;
aud[34564]=16'h3cff;
aud[34565]=16'h3d05;
aud[34566]=16'h3d0c;
aud[34567]=16'h3d12;
aud[34568]=16'h3d19;
aud[34569]=16'h3d1f;
aud[34570]=16'h3d25;
aud[34571]=16'h3d2c;
aud[34572]=16'h3d32;
aud[34573]=16'h3d38;
aud[34574]=16'h3d3f;
aud[34575]=16'h3d45;
aud[34576]=16'h3d4b;
aud[34577]=16'h3d51;
aud[34578]=16'h3d57;
aud[34579]=16'h3d5d;
aud[34580]=16'h3d63;
aud[34581]=16'h3d69;
aud[34582]=16'h3d6f;
aud[34583]=16'h3d75;
aud[34584]=16'h3d7b;
aud[34585]=16'h3d81;
aud[34586]=16'h3d87;
aud[34587]=16'h3d8d;
aud[34588]=16'h3d93;
aud[34589]=16'h3d99;
aud[34590]=16'h3d9f;
aud[34591]=16'h3da4;
aud[34592]=16'h3daa;
aud[34593]=16'h3db0;
aud[34594]=16'h3db6;
aud[34595]=16'h3dbb;
aud[34596]=16'h3dc1;
aud[34597]=16'h3dc7;
aud[34598]=16'h3dcc;
aud[34599]=16'h3dd2;
aud[34600]=16'h3dd7;
aud[34601]=16'h3ddd;
aud[34602]=16'h3de2;
aud[34603]=16'h3de8;
aud[34604]=16'h3ded;
aud[34605]=16'h3df3;
aud[34606]=16'h3df8;
aud[34607]=16'h3dfd;
aud[34608]=16'h3e03;
aud[34609]=16'h3e08;
aud[34610]=16'h3e0d;
aud[34611]=16'h3e12;
aud[34612]=16'h3e18;
aud[34613]=16'h3e1d;
aud[34614]=16'h3e22;
aud[34615]=16'h3e27;
aud[34616]=16'h3e2c;
aud[34617]=16'h3e31;
aud[34618]=16'h3e36;
aud[34619]=16'h3e3b;
aud[34620]=16'h3e40;
aud[34621]=16'h3e45;
aud[34622]=16'h3e4a;
aud[34623]=16'h3e4f;
aud[34624]=16'h3e54;
aud[34625]=16'h3e59;
aud[34626]=16'h3e5e;
aud[34627]=16'h3e62;
aud[34628]=16'h3e67;
aud[34629]=16'h3e6c;
aud[34630]=16'h3e71;
aud[34631]=16'h3e75;
aud[34632]=16'h3e7a;
aud[34633]=16'h3e7f;
aud[34634]=16'h3e83;
aud[34635]=16'h3e88;
aud[34636]=16'h3e8c;
aud[34637]=16'h3e91;
aud[34638]=16'h3e95;
aud[34639]=16'h3e9a;
aud[34640]=16'h3e9e;
aud[34641]=16'h3ea3;
aud[34642]=16'h3ea7;
aud[34643]=16'h3eac;
aud[34644]=16'h3eb0;
aud[34645]=16'h3eb4;
aud[34646]=16'h3eb9;
aud[34647]=16'h3ebd;
aud[34648]=16'h3ec1;
aud[34649]=16'h3ec5;
aud[34650]=16'h3ec9;
aud[34651]=16'h3ecd;
aud[34652]=16'h3ed2;
aud[34653]=16'h3ed6;
aud[34654]=16'h3eda;
aud[34655]=16'h3ede;
aud[34656]=16'h3ee2;
aud[34657]=16'h3ee6;
aud[34658]=16'h3eea;
aud[34659]=16'h3eee;
aud[34660]=16'h3ef2;
aud[34661]=16'h3ef5;
aud[34662]=16'h3ef9;
aud[34663]=16'h3efd;
aud[34664]=16'h3f01;
aud[34665]=16'h3f05;
aud[34666]=16'h3f08;
aud[34667]=16'h3f0c;
aud[34668]=16'h3f10;
aud[34669]=16'h3f13;
aud[34670]=16'h3f17;
aud[34671]=16'h3f1b;
aud[34672]=16'h3f1e;
aud[34673]=16'h3f22;
aud[34674]=16'h3f25;
aud[34675]=16'h3f29;
aud[34676]=16'h3f2c;
aud[34677]=16'h3f30;
aud[34678]=16'h3f33;
aud[34679]=16'h3f36;
aud[34680]=16'h3f3a;
aud[34681]=16'h3f3d;
aud[34682]=16'h3f40;
aud[34683]=16'h3f43;
aud[34684]=16'h3f47;
aud[34685]=16'h3f4a;
aud[34686]=16'h3f4d;
aud[34687]=16'h3f50;
aud[34688]=16'h3f53;
aud[34689]=16'h3f56;
aud[34690]=16'h3f5a;
aud[34691]=16'h3f5d;
aud[34692]=16'h3f60;
aud[34693]=16'h3f63;
aud[34694]=16'h3f65;
aud[34695]=16'h3f68;
aud[34696]=16'h3f6b;
aud[34697]=16'h3f6e;
aud[34698]=16'h3f71;
aud[34699]=16'h3f74;
aud[34700]=16'h3f77;
aud[34701]=16'h3f79;
aud[34702]=16'h3f7c;
aud[34703]=16'h3f7f;
aud[34704]=16'h3f81;
aud[34705]=16'h3f84;
aud[34706]=16'h3f87;
aud[34707]=16'h3f89;
aud[34708]=16'h3f8c;
aud[34709]=16'h3f8e;
aud[34710]=16'h3f91;
aud[34711]=16'h3f93;
aud[34712]=16'h3f96;
aud[34713]=16'h3f98;
aud[34714]=16'h3f9b;
aud[34715]=16'h3f9d;
aud[34716]=16'h3f9f;
aud[34717]=16'h3fa2;
aud[34718]=16'h3fa4;
aud[34719]=16'h3fa6;
aud[34720]=16'h3fa8;
aud[34721]=16'h3fab;
aud[34722]=16'h3fad;
aud[34723]=16'h3faf;
aud[34724]=16'h3fb1;
aud[34725]=16'h3fb3;
aud[34726]=16'h3fb5;
aud[34727]=16'h3fb7;
aud[34728]=16'h3fb9;
aud[34729]=16'h3fbb;
aud[34730]=16'h3fbd;
aud[34731]=16'h3fbf;
aud[34732]=16'h3fc1;
aud[34733]=16'h3fc3;
aud[34734]=16'h3fc5;
aud[34735]=16'h3fc7;
aud[34736]=16'h3fc8;
aud[34737]=16'h3fca;
aud[34738]=16'h3fcc;
aud[34739]=16'h3fcd;
aud[34740]=16'h3fcf;
aud[34741]=16'h3fd1;
aud[34742]=16'h3fd2;
aud[34743]=16'h3fd4;
aud[34744]=16'h3fd6;
aud[34745]=16'h3fd7;
aud[34746]=16'h3fd9;
aud[34747]=16'h3fda;
aud[34748]=16'h3fdc;
aud[34749]=16'h3fdd;
aud[34750]=16'h3fde;
aud[34751]=16'h3fe0;
aud[34752]=16'h3fe1;
aud[34753]=16'h3fe2;
aud[34754]=16'h3fe4;
aud[34755]=16'h3fe5;
aud[34756]=16'h3fe6;
aud[34757]=16'h3fe7;
aud[34758]=16'h3fe8;
aud[34759]=16'h3fea;
aud[34760]=16'h3feb;
aud[34761]=16'h3fec;
aud[34762]=16'h3fed;
aud[34763]=16'h3fee;
aud[34764]=16'h3fef;
aud[34765]=16'h3ff0;
aud[34766]=16'h3ff1;
aud[34767]=16'h3ff2;
aud[34768]=16'h3ff3;
aud[34769]=16'h3ff3;
aud[34770]=16'h3ff4;
aud[34771]=16'h3ff5;
aud[34772]=16'h3ff6;
aud[34773]=16'h3ff7;
aud[34774]=16'h3ff7;
aud[34775]=16'h3ff8;
aud[34776]=16'h3ff9;
aud[34777]=16'h3ff9;
aud[34778]=16'h3ffa;
aud[34779]=16'h3ffa;
aud[34780]=16'h3ffb;
aud[34781]=16'h3ffb;
aud[34782]=16'h3ffc;
aud[34783]=16'h3ffc;
aud[34784]=16'h3ffd;
aud[34785]=16'h3ffd;
aud[34786]=16'h3ffe;
aud[34787]=16'h3ffe;
aud[34788]=16'h3ffe;
aud[34789]=16'h3fff;
aud[34790]=16'h3fff;
aud[34791]=16'h3fff;
aud[34792]=16'h3fff;
aud[34793]=16'h3fff;
aud[34794]=16'h4000;
aud[34795]=16'h4000;
aud[34796]=16'h4000;
aud[34797]=16'h4000;
aud[34798]=16'h4000;
aud[34799]=16'h4000;
aud[34800]=16'h4000;
aud[34801]=16'h4000;
aud[34802]=16'h4000;
aud[34803]=16'h4000;
aud[34804]=16'h4000;
aud[34805]=16'h3fff;
aud[34806]=16'h3fff;
aud[34807]=16'h3fff;
aud[34808]=16'h3fff;
aud[34809]=16'h3fff;
aud[34810]=16'h3ffe;
aud[34811]=16'h3ffe;
aud[34812]=16'h3ffe;
aud[34813]=16'h3ffd;
aud[34814]=16'h3ffd;
aud[34815]=16'h3ffc;
aud[34816]=16'h3ffc;
aud[34817]=16'h3ffb;
aud[34818]=16'h3ffb;
aud[34819]=16'h3ffa;
aud[34820]=16'h3ffa;
aud[34821]=16'h3ff9;
aud[34822]=16'h3ff9;
aud[34823]=16'h3ff8;
aud[34824]=16'h3ff7;
aud[34825]=16'h3ff7;
aud[34826]=16'h3ff6;
aud[34827]=16'h3ff5;
aud[34828]=16'h3ff4;
aud[34829]=16'h3ff3;
aud[34830]=16'h3ff3;
aud[34831]=16'h3ff2;
aud[34832]=16'h3ff1;
aud[34833]=16'h3ff0;
aud[34834]=16'h3fef;
aud[34835]=16'h3fee;
aud[34836]=16'h3fed;
aud[34837]=16'h3fec;
aud[34838]=16'h3feb;
aud[34839]=16'h3fea;
aud[34840]=16'h3fe8;
aud[34841]=16'h3fe7;
aud[34842]=16'h3fe6;
aud[34843]=16'h3fe5;
aud[34844]=16'h3fe4;
aud[34845]=16'h3fe2;
aud[34846]=16'h3fe1;
aud[34847]=16'h3fe0;
aud[34848]=16'h3fde;
aud[34849]=16'h3fdd;
aud[34850]=16'h3fdc;
aud[34851]=16'h3fda;
aud[34852]=16'h3fd9;
aud[34853]=16'h3fd7;
aud[34854]=16'h3fd6;
aud[34855]=16'h3fd4;
aud[34856]=16'h3fd2;
aud[34857]=16'h3fd1;
aud[34858]=16'h3fcf;
aud[34859]=16'h3fcd;
aud[34860]=16'h3fcc;
aud[34861]=16'h3fca;
aud[34862]=16'h3fc8;
aud[34863]=16'h3fc7;
aud[34864]=16'h3fc5;
aud[34865]=16'h3fc3;
aud[34866]=16'h3fc1;
aud[34867]=16'h3fbf;
aud[34868]=16'h3fbd;
aud[34869]=16'h3fbb;
aud[34870]=16'h3fb9;
aud[34871]=16'h3fb7;
aud[34872]=16'h3fb5;
aud[34873]=16'h3fb3;
aud[34874]=16'h3fb1;
aud[34875]=16'h3faf;
aud[34876]=16'h3fad;
aud[34877]=16'h3fab;
aud[34878]=16'h3fa8;
aud[34879]=16'h3fa6;
aud[34880]=16'h3fa4;
aud[34881]=16'h3fa2;
aud[34882]=16'h3f9f;
aud[34883]=16'h3f9d;
aud[34884]=16'h3f9b;
aud[34885]=16'h3f98;
aud[34886]=16'h3f96;
aud[34887]=16'h3f93;
aud[34888]=16'h3f91;
aud[34889]=16'h3f8e;
aud[34890]=16'h3f8c;
aud[34891]=16'h3f89;
aud[34892]=16'h3f87;
aud[34893]=16'h3f84;
aud[34894]=16'h3f81;
aud[34895]=16'h3f7f;
aud[34896]=16'h3f7c;
aud[34897]=16'h3f79;
aud[34898]=16'h3f77;
aud[34899]=16'h3f74;
aud[34900]=16'h3f71;
aud[34901]=16'h3f6e;
aud[34902]=16'h3f6b;
aud[34903]=16'h3f68;
aud[34904]=16'h3f65;
aud[34905]=16'h3f63;
aud[34906]=16'h3f60;
aud[34907]=16'h3f5d;
aud[34908]=16'h3f5a;
aud[34909]=16'h3f56;
aud[34910]=16'h3f53;
aud[34911]=16'h3f50;
aud[34912]=16'h3f4d;
aud[34913]=16'h3f4a;
aud[34914]=16'h3f47;
aud[34915]=16'h3f43;
aud[34916]=16'h3f40;
aud[34917]=16'h3f3d;
aud[34918]=16'h3f3a;
aud[34919]=16'h3f36;
aud[34920]=16'h3f33;
aud[34921]=16'h3f30;
aud[34922]=16'h3f2c;
aud[34923]=16'h3f29;
aud[34924]=16'h3f25;
aud[34925]=16'h3f22;
aud[34926]=16'h3f1e;
aud[34927]=16'h3f1b;
aud[34928]=16'h3f17;
aud[34929]=16'h3f13;
aud[34930]=16'h3f10;
aud[34931]=16'h3f0c;
aud[34932]=16'h3f08;
aud[34933]=16'h3f05;
aud[34934]=16'h3f01;
aud[34935]=16'h3efd;
aud[34936]=16'h3ef9;
aud[34937]=16'h3ef5;
aud[34938]=16'h3ef2;
aud[34939]=16'h3eee;
aud[34940]=16'h3eea;
aud[34941]=16'h3ee6;
aud[34942]=16'h3ee2;
aud[34943]=16'h3ede;
aud[34944]=16'h3eda;
aud[34945]=16'h3ed6;
aud[34946]=16'h3ed2;
aud[34947]=16'h3ecd;
aud[34948]=16'h3ec9;
aud[34949]=16'h3ec5;
aud[34950]=16'h3ec1;
aud[34951]=16'h3ebd;
aud[34952]=16'h3eb9;
aud[34953]=16'h3eb4;
aud[34954]=16'h3eb0;
aud[34955]=16'h3eac;
aud[34956]=16'h3ea7;
aud[34957]=16'h3ea3;
aud[34958]=16'h3e9e;
aud[34959]=16'h3e9a;
aud[34960]=16'h3e95;
aud[34961]=16'h3e91;
aud[34962]=16'h3e8c;
aud[34963]=16'h3e88;
aud[34964]=16'h3e83;
aud[34965]=16'h3e7f;
aud[34966]=16'h3e7a;
aud[34967]=16'h3e75;
aud[34968]=16'h3e71;
aud[34969]=16'h3e6c;
aud[34970]=16'h3e67;
aud[34971]=16'h3e62;
aud[34972]=16'h3e5e;
aud[34973]=16'h3e59;
aud[34974]=16'h3e54;
aud[34975]=16'h3e4f;
aud[34976]=16'h3e4a;
aud[34977]=16'h3e45;
aud[34978]=16'h3e40;
aud[34979]=16'h3e3b;
aud[34980]=16'h3e36;
aud[34981]=16'h3e31;
aud[34982]=16'h3e2c;
aud[34983]=16'h3e27;
aud[34984]=16'h3e22;
aud[34985]=16'h3e1d;
aud[34986]=16'h3e18;
aud[34987]=16'h3e12;
aud[34988]=16'h3e0d;
aud[34989]=16'h3e08;
aud[34990]=16'h3e03;
aud[34991]=16'h3dfd;
aud[34992]=16'h3df8;
aud[34993]=16'h3df3;
aud[34994]=16'h3ded;
aud[34995]=16'h3de8;
aud[34996]=16'h3de2;
aud[34997]=16'h3ddd;
aud[34998]=16'h3dd7;
aud[34999]=16'h3dd2;
aud[35000]=16'h3dcc;
aud[35001]=16'h3dc7;
aud[35002]=16'h3dc1;
aud[35003]=16'h3dbb;
aud[35004]=16'h3db6;
aud[35005]=16'h3db0;
aud[35006]=16'h3daa;
aud[35007]=16'h3da4;
aud[35008]=16'h3d9f;
aud[35009]=16'h3d99;
aud[35010]=16'h3d93;
aud[35011]=16'h3d8d;
aud[35012]=16'h3d87;
aud[35013]=16'h3d81;
aud[35014]=16'h3d7b;
aud[35015]=16'h3d75;
aud[35016]=16'h3d6f;
aud[35017]=16'h3d69;
aud[35018]=16'h3d63;
aud[35019]=16'h3d5d;
aud[35020]=16'h3d57;
aud[35021]=16'h3d51;
aud[35022]=16'h3d4b;
aud[35023]=16'h3d45;
aud[35024]=16'h3d3f;
aud[35025]=16'h3d38;
aud[35026]=16'h3d32;
aud[35027]=16'h3d2c;
aud[35028]=16'h3d25;
aud[35029]=16'h3d1f;
aud[35030]=16'h3d19;
aud[35031]=16'h3d12;
aud[35032]=16'h3d0c;
aud[35033]=16'h3d05;
aud[35034]=16'h3cff;
aud[35035]=16'h3cf8;
aud[35036]=16'h3cf2;
aud[35037]=16'h3ceb;
aud[35038]=16'h3ce5;
aud[35039]=16'h3cde;
aud[35040]=16'h3cd7;
aud[35041]=16'h3cd1;
aud[35042]=16'h3cca;
aud[35043]=16'h3cc3;
aud[35044]=16'h3cbd;
aud[35045]=16'h3cb6;
aud[35046]=16'h3caf;
aud[35047]=16'h3ca8;
aud[35048]=16'h3ca1;
aud[35049]=16'h3c9b;
aud[35050]=16'h3c94;
aud[35051]=16'h3c8d;
aud[35052]=16'h3c86;
aud[35053]=16'h3c7f;
aud[35054]=16'h3c78;
aud[35055]=16'h3c71;
aud[35056]=16'h3c6a;
aud[35057]=16'h3c63;
aud[35058]=16'h3c5b;
aud[35059]=16'h3c54;
aud[35060]=16'h3c4d;
aud[35061]=16'h3c46;
aud[35062]=16'h3c3f;
aud[35063]=16'h3c37;
aud[35064]=16'h3c30;
aud[35065]=16'h3c29;
aud[35066]=16'h3c21;
aud[35067]=16'h3c1a;
aud[35068]=16'h3c13;
aud[35069]=16'h3c0b;
aud[35070]=16'h3c04;
aud[35071]=16'h3bfc;
aud[35072]=16'h3bf5;
aud[35073]=16'h3bed;
aud[35074]=16'h3be6;
aud[35075]=16'h3bde;
aud[35076]=16'h3bd7;
aud[35077]=16'h3bcf;
aud[35078]=16'h3bc7;
aud[35079]=16'h3bc0;
aud[35080]=16'h3bb8;
aud[35081]=16'h3bb0;
aud[35082]=16'h3ba9;
aud[35083]=16'h3ba1;
aud[35084]=16'h3b99;
aud[35085]=16'h3b91;
aud[35086]=16'h3b89;
aud[35087]=16'h3b81;
aud[35088]=16'h3b7a;
aud[35089]=16'h3b72;
aud[35090]=16'h3b6a;
aud[35091]=16'h3b62;
aud[35092]=16'h3b5a;
aud[35093]=16'h3b52;
aud[35094]=16'h3b4a;
aud[35095]=16'h3b41;
aud[35096]=16'h3b39;
aud[35097]=16'h3b31;
aud[35098]=16'h3b29;
aud[35099]=16'h3b21;
aud[35100]=16'h3b19;
aud[35101]=16'h3b10;
aud[35102]=16'h3b08;
aud[35103]=16'h3b00;
aud[35104]=16'h3af7;
aud[35105]=16'h3aef;
aud[35106]=16'h3ae7;
aud[35107]=16'h3ade;
aud[35108]=16'h3ad6;
aud[35109]=16'h3acd;
aud[35110]=16'h3ac5;
aud[35111]=16'h3abc;
aud[35112]=16'h3ab4;
aud[35113]=16'h3aab;
aud[35114]=16'h3aa3;
aud[35115]=16'h3a9a;
aud[35116]=16'h3a92;
aud[35117]=16'h3a89;
aud[35118]=16'h3a80;
aud[35119]=16'h3a78;
aud[35120]=16'h3a6f;
aud[35121]=16'h3a66;
aud[35122]=16'h3a5d;
aud[35123]=16'h3a54;
aud[35124]=16'h3a4c;
aud[35125]=16'h3a43;
aud[35126]=16'h3a3a;
aud[35127]=16'h3a31;
aud[35128]=16'h3a28;
aud[35129]=16'h3a1f;
aud[35130]=16'h3a16;
aud[35131]=16'h3a0d;
aud[35132]=16'h3a04;
aud[35133]=16'h39fb;
aud[35134]=16'h39f2;
aud[35135]=16'h39e9;
aud[35136]=16'h39e0;
aud[35137]=16'h39d6;
aud[35138]=16'h39cd;
aud[35139]=16'h39c4;
aud[35140]=16'h39bb;
aud[35141]=16'h39b1;
aud[35142]=16'h39a8;
aud[35143]=16'h399f;
aud[35144]=16'h3995;
aud[35145]=16'h398c;
aud[35146]=16'h3983;
aud[35147]=16'h3979;
aud[35148]=16'h3970;
aud[35149]=16'h3966;
aud[35150]=16'h395d;
aud[35151]=16'h3953;
aud[35152]=16'h394a;
aud[35153]=16'h3940;
aud[35154]=16'h3937;
aud[35155]=16'h392d;
aud[35156]=16'h3923;
aud[35157]=16'h391a;
aud[35158]=16'h3910;
aud[35159]=16'h3906;
aud[35160]=16'h38fd;
aud[35161]=16'h38f3;
aud[35162]=16'h38e9;
aud[35163]=16'h38df;
aud[35164]=16'h38d5;
aud[35165]=16'h38cb;
aud[35166]=16'h38c1;
aud[35167]=16'h38b8;
aud[35168]=16'h38ae;
aud[35169]=16'h38a4;
aud[35170]=16'h389a;
aud[35171]=16'h3890;
aud[35172]=16'h3886;
aud[35173]=16'h387b;
aud[35174]=16'h3871;
aud[35175]=16'h3867;
aud[35176]=16'h385d;
aud[35177]=16'h3853;
aud[35178]=16'h3849;
aud[35179]=16'h383f;
aud[35180]=16'h3834;
aud[35181]=16'h382a;
aud[35182]=16'h3820;
aud[35183]=16'h3815;
aud[35184]=16'h380b;
aud[35185]=16'h3801;
aud[35186]=16'h37f6;
aud[35187]=16'h37ec;
aud[35188]=16'h37e1;
aud[35189]=16'h37d7;
aud[35190]=16'h37cc;
aud[35191]=16'h37c2;
aud[35192]=16'h37b7;
aud[35193]=16'h37ad;
aud[35194]=16'h37a2;
aud[35195]=16'h3798;
aud[35196]=16'h378d;
aud[35197]=16'h3782;
aud[35198]=16'h3778;
aud[35199]=16'h376d;
aud[35200]=16'h3762;
aud[35201]=16'h3757;
aud[35202]=16'h374d;
aud[35203]=16'h3742;
aud[35204]=16'h3737;
aud[35205]=16'h372c;
aud[35206]=16'h3721;
aud[35207]=16'h3716;
aud[35208]=16'h370b;
aud[35209]=16'h3701;
aud[35210]=16'h36f6;
aud[35211]=16'h36eb;
aud[35212]=16'h36e0;
aud[35213]=16'h36d4;
aud[35214]=16'h36c9;
aud[35215]=16'h36be;
aud[35216]=16'h36b3;
aud[35217]=16'h36a8;
aud[35218]=16'h369d;
aud[35219]=16'h3692;
aud[35220]=16'h3686;
aud[35221]=16'h367b;
aud[35222]=16'h3670;
aud[35223]=16'h3665;
aud[35224]=16'h3659;
aud[35225]=16'h364e;
aud[35226]=16'h3643;
aud[35227]=16'h3637;
aud[35228]=16'h362c;
aud[35229]=16'h3620;
aud[35230]=16'h3615;
aud[35231]=16'h3609;
aud[35232]=16'h35fe;
aud[35233]=16'h35f2;
aud[35234]=16'h35e7;
aud[35235]=16'h35db;
aud[35236]=16'h35d0;
aud[35237]=16'h35c4;
aud[35238]=16'h35b8;
aud[35239]=16'h35ad;
aud[35240]=16'h35a1;
aud[35241]=16'h3595;
aud[35242]=16'h358a;
aud[35243]=16'h357e;
aud[35244]=16'h3572;
aud[35245]=16'h3566;
aud[35246]=16'h355a;
aud[35247]=16'h354f;
aud[35248]=16'h3543;
aud[35249]=16'h3537;
aud[35250]=16'h352b;
aud[35251]=16'h351f;
aud[35252]=16'h3513;
aud[35253]=16'h3507;
aud[35254]=16'h34fb;
aud[35255]=16'h34ef;
aud[35256]=16'h34e3;
aud[35257]=16'h34d7;
aud[35258]=16'h34cb;
aud[35259]=16'h34be;
aud[35260]=16'h34b2;
aud[35261]=16'h34a6;
aud[35262]=16'h349a;
aud[35263]=16'h348e;
aud[35264]=16'h3481;
aud[35265]=16'h3475;
aud[35266]=16'h3469;
aud[35267]=16'h345d;
aud[35268]=16'h3450;
aud[35269]=16'h3444;
aud[35270]=16'h3437;
aud[35271]=16'h342b;
aud[35272]=16'h341f;
aud[35273]=16'h3412;
aud[35274]=16'h3406;
aud[35275]=16'h33f9;
aud[35276]=16'h33ed;
aud[35277]=16'h33e0;
aud[35278]=16'h33d4;
aud[35279]=16'h33c7;
aud[35280]=16'h33ba;
aud[35281]=16'h33ae;
aud[35282]=16'h33a1;
aud[35283]=16'h3394;
aud[35284]=16'h3388;
aud[35285]=16'h337b;
aud[35286]=16'h336e;
aud[35287]=16'h3361;
aud[35288]=16'h3355;
aud[35289]=16'h3348;
aud[35290]=16'h333b;
aud[35291]=16'h332e;
aud[35292]=16'h3321;
aud[35293]=16'h3314;
aud[35294]=16'h3307;
aud[35295]=16'h32fa;
aud[35296]=16'h32ed;
aud[35297]=16'h32e0;
aud[35298]=16'h32d3;
aud[35299]=16'h32c6;
aud[35300]=16'h32b9;
aud[35301]=16'h32ac;
aud[35302]=16'h329f;
aud[35303]=16'h3292;
aud[35304]=16'h3285;
aud[35305]=16'h3278;
aud[35306]=16'h326a;
aud[35307]=16'h325d;
aud[35308]=16'h3250;
aud[35309]=16'h3243;
aud[35310]=16'h3235;
aud[35311]=16'h3228;
aud[35312]=16'h321b;
aud[35313]=16'h320d;
aud[35314]=16'h3200;
aud[35315]=16'h31f3;
aud[35316]=16'h31e5;
aud[35317]=16'h31d8;
aud[35318]=16'h31ca;
aud[35319]=16'h31bd;
aud[35320]=16'h31af;
aud[35321]=16'h31a2;
aud[35322]=16'h3194;
aud[35323]=16'h3187;
aud[35324]=16'h3179;
aud[35325]=16'h316b;
aud[35326]=16'h315e;
aud[35327]=16'h3150;
aud[35328]=16'h3142;
aud[35329]=16'h3135;
aud[35330]=16'h3127;
aud[35331]=16'h3119;
aud[35332]=16'h310b;
aud[35333]=16'h30fe;
aud[35334]=16'h30f0;
aud[35335]=16'h30e2;
aud[35336]=16'h30d4;
aud[35337]=16'h30c6;
aud[35338]=16'h30b8;
aud[35339]=16'h30aa;
aud[35340]=16'h309d;
aud[35341]=16'h308f;
aud[35342]=16'h3081;
aud[35343]=16'h3073;
aud[35344]=16'h3065;
aud[35345]=16'h3057;
aud[35346]=16'h3048;
aud[35347]=16'h303a;
aud[35348]=16'h302c;
aud[35349]=16'h301e;
aud[35350]=16'h3010;
aud[35351]=16'h3002;
aud[35352]=16'h2ff4;
aud[35353]=16'h2fe5;
aud[35354]=16'h2fd7;
aud[35355]=16'h2fc9;
aud[35356]=16'h2fbb;
aud[35357]=16'h2fac;
aud[35358]=16'h2f9e;
aud[35359]=16'h2f90;
aud[35360]=16'h2f81;
aud[35361]=16'h2f73;
aud[35362]=16'h2f65;
aud[35363]=16'h2f56;
aud[35364]=16'h2f48;
aud[35365]=16'h2f39;
aud[35366]=16'h2f2b;
aud[35367]=16'h2f1c;
aud[35368]=16'h2f0e;
aud[35369]=16'h2eff;
aud[35370]=16'h2ef1;
aud[35371]=16'h2ee2;
aud[35372]=16'h2ed3;
aud[35373]=16'h2ec5;
aud[35374]=16'h2eb6;
aud[35375]=16'h2ea7;
aud[35376]=16'h2e99;
aud[35377]=16'h2e8a;
aud[35378]=16'h2e7b;
aud[35379]=16'h2e6d;
aud[35380]=16'h2e5e;
aud[35381]=16'h2e4f;
aud[35382]=16'h2e40;
aud[35383]=16'h2e31;
aud[35384]=16'h2e22;
aud[35385]=16'h2e14;
aud[35386]=16'h2e05;
aud[35387]=16'h2df6;
aud[35388]=16'h2de7;
aud[35389]=16'h2dd8;
aud[35390]=16'h2dc9;
aud[35391]=16'h2dba;
aud[35392]=16'h2dab;
aud[35393]=16'h2d9c;
aud[35394]=16'h2d8d;
aud[35395]=16'h2d7e;
aud[35396]=16'h2d6f;
aud[35397]=16'h2d60;
aud[35398]=16'h2d50;
aud[35399]=16'h2d41;
aud[35400]=16'h2d32;
aud[35401]=16'h2d23;
aud[35402]=16'h2d14;
aud[35403]=16'h2d04;
aud[35404]=16'h2cf5;
aud[35405]=16'h2ce6;
aud[35406]=16'h2cd7;
aud[35407]=16'h2cc7;
aud[35408]=16'h2cb8;
aud[35409]=16'h2ca9;
aud[35410]=16'h2c99;
aud[35411]=16'h2c8a;
aud[35412]=16'h2c7a;
aud[35413]=16'h2c6b;
aud[35414]=16'h2c5c;
aud[35415]=16'h2c4c;
aud[35416]=16'h2c3d;
aud[35417]=16'h2c2d;
aud[35418]=16'h2c1e;
aud[35419]=16'h2c0e;
aud[35420]=16'h2bfe;
aud[35421]=16'h2bef;
aud[35422]=16'h2bdf;
aud[35423]=16'h2bd0;
aud[35424]=16'h2bc0;
aud[35425]=16'h2bb0;
aud[35426]=16'h2ba1;
aud[35427]=16'h2b91;
aud[35428]=16'h2b81;
aud[35429]=16'h2b71;
aud[35430]=16'h2b62;
aud[35431]=16'h2b52;
aud[35432]=16'h2b42;
aud[35433]=16'h2b32;
aud[35434]=16'h2b22;
aud[35435]=16'h2b13;
aud[35436]=16'h2b03;
aud[35437]=16'h2af3;
aud[35438]=16'h2ae3;
aud[35439]=16'h2ad3;
aud[35440]=16'h2ac3;
aud[35441]=16'h2ab3;
aud[35442]=16'h2aa3;
aud[35443]=16'h2a93;
aud[35444]=16'h2a83;
aud[35445]=16'h2a73;
aud[35446]=16'h2a63;
aud[35447]=16'h2a53;
aud[35448]=16'h2a43;
aud[35449]=16'h2a33;
aud[35450]=16'h2a23;
aud[35451]=16'h2a12;
aud[35452]=16'h2a02;
aud[35453]=16'h29f2;
aud[35454]=16'h29e2;
aud[35455]=16'h29d2;
aud[35456]=16'h29c1;
aud[35457]=16'h29b1;
aud[35458]=16'h29a1;
aud[35459]=16'h2991;
aud[35460]=16'h2980;
aud[35461]=16'h2970;
aud[35462]=16'h2960;
aud[35463]=16'h294f;
aud[35464]=16'h293f;
aud[35465]=16'h292e;
aud[35466]=16'h291e;
aud[35467]=16'h290e;
aud[35468]=16'h28fd;
aud[35469]=16'h28ed;
aud[35470]=16'h28dc;
aud[35471]=16'h28cc;
aud[35472]=16'h28bb;
aud[35473]=16'h28aa;
aud[35474]=16'h289a;
aud[35475]=16'h2889;
aud[35476]=16'h2879;
aud[35477]=16'h2868;
aud[35478]=16'h2857;
aud[35479]=16'h2847;
aud[35480]=16'h2836;
aud[35481]=16'h2825;
aud[35482]=16'h2815;
aud[35483]=16'h2804;
aud[35484]=16'h27f3;
aud[35485]=16'h27e2;
aud[35486]=16'h27d2;
aud[35487]=16'h27c1;
aud[35488]=16'h27b0;
aud[35489]=16'h279f;
aud[35490]=16'h278e;
aud[35491]=16'h277e;
aud[35492]=16'h276d;
aud[35493]=16'h275c;
aud[35494]=16'h274b;
aud[35495]=16'h273a;
aud[35496]=16'h2729;
aud[35497]=16'h2718;
aud[35498]=16'h2707;
aud[35499]=16'h26f6;
aud[35500]=16'h26e5;
aud[35501]=16'h26d4;
aud[35502]=16'h26c3;
aud[35503]=16'h26b2;
aud[35504]=16'h26a1;
aud[35505]=16'h2690;
aud[35506]=16'h267e;
aud[35507]=16'h266d;
aud[35508]=16'h265c;
aud[35509]=16'h264b;
aud[35510]=16'h263a;
aud[35511]=16'h2629;
aud[35512]=16'h2617;
aud[35513]=16'h2606;
aud[35514]=16'h25f5;
aud[35515]=16'h25e4;
aud[35516]=16'h25d2;
aud[35517]=16'h25c1;
aud[35518]=16'h25b0;
aud[35519]=16'h259e;
aud[35520]=16'h258d;
aud[35521]=16'h257c;
aud[35522]=16'h256a;
aud[35523]=16'h2559;
aud[35524]=16'h2547;
aud[35525]=16'h2536;
aud[35526]=16'h2524;
aud[35527]=16'h2513;
aud[35528]=16'h2501;
aud[35529]=16'h24f0;
aud[35530]=16'h24de;
aud[35531]=16'h24cd;
aud[35532]=16'h24bb;
aud[35533]=16'h24aa;
aud[35534]=16'h2498;
aud[35535]=16'h2487;
aud[35536]=16'h2475;
aud[35537]=16'h2463;
aud[35538]=16'h2452;
aud[35539]=16'h2440;
aud[35540]=16'h242e;
aud[35541]=16'h241d;
aud[35542]=16'h240b;
aud[35543]=16'h23f9;
aud[35544]=16'h23e7;
aud[35545]=16'h23d6;
aud[35546]=16'h23c4;
aud[35547]=16'h23b2;
aud[35548]=16'h23a0;
aud[35549]=16'h238e;
aud[35550]=16'h237d;
aud[35551]=16'h236b;
aud[35552]=16'h2359;
aud[35553]=16'h2347;
aud[35554]=16'h2335;
aud[35555]=16'h2323;
aud[35556]=16'h2311;
aud[35557]=16'h22ff;
aud[35558]=16'h22ed;
aud[35559]=16'h22db;
aud[35560]=16'h22c9;
aud[35561]=16'h22b7;
aud[35562]=16'h22a5;
aud[35563]=16'h2293;
aud[35564]=16'h2281;
aud[35565]=16'h226f;
aud[35566]=16'h225d;
aud[35567]=16'h224b;
aud[35568]=16'h2239;
aud[35569]=16'h2227;
aud[35570]=16'h2215;
aud[35571]=16'h2202;
aud[35572]=16'h21f0;
aud[35573]=16'h21de;
aud[35574]=16'h21cc;
aud[35575]=16'h21ba;
aud[35576]=16'h21a7;
aud[35577]=16'h2195;
aud[35578]=16'h2183;
aud[35579]=16'h2171;
aud[35580]=16'h215e;
aud[35581]=16'h214c;
aud[35582]=16'h213a;
aud[35583]=16'h2127;
aud[35584]=16'h2115;
aud[35585]=16'h2103;
aud[35586]=16'h20f0;
aud[35587]=16'h20de;
aud[35588]=16'h20cb;
aud[35589]=16'h20b9;
aud[35590]=16'h20a7;
aud[35591]=16'h2094;
aud[35592]=16'h2082;
aud[35593]=16'h206f;
aud[35594]=16'h205d;
aud[35595]=16'h204a;
aud[35596]=16'h2038;
aud[35597]=16'h2025;
aud[35598]=16'h2013;
aud[35599]=16'h2000;
aud[35600]=16'h1fed;
aud[35601]=16'h1fdb;
aud[35602]=16'h1fc8;
aud[35603]=16'h1fb6;
aud[35604]=16'h1fa3;
aud[35605]=16'h1f90;
aud[35606]=16'h1f7e;
aud[35607]=16'h1f6b;
aud[35608]=16'h1f58;
aud[35609]=16'h1f46;
aud[35610]=16'h1f33;
aud[35611]=16'h1f20;
aud[35612]=16'h1f0d;
aud[35613]=16'h1efb;
aud[35614]=16'h1ee8;
aud[35615]=16'h1ed5;
aud[35616]=16'h1ec2;
aud[35617]=16'h1eaf;
aud[35618]=16'h1e9d;
aud[35619]=16'h1e8a;
aud[35620]=16'h1e77;
aud[35621]=16'h1e64;
aud[35622]=16'h1e51;
aud[35623]=16'h1e3e;
aud[35624]=16'h1e2b;
aud[35625]=16'h1e18;
aud[35626]=16'h1e06;
aud[35627]=16'h1df3;
aud[35628]=16'h1de0;
aud[35629]=16'h1dcd;
aud[35630]=16'h1dba;
aud[35631]=16'h1da7;
aud[35632]=16'h1d94;
aud[35633]=16'h1d81;
aud[35634]=16'h1d6e;
aud[35635]=16'h1d5b;
aud[35636]=16'h1d47;
aud[35637]=16'h1d34;
aud[35638]=16'h1d21;
aud[35639]=16'h1d0e;
aud[35640]=16'h1cfb;
aud[35641]=16'h1ce8;
aud[35642]=16'h1cd5;
aud[35643]=16'h1cc2;
aud[35644]=16'h1cae;
aud[35645]=16'h1c9b;
aud[35646]=16'h1c88;
aud[35647]=16'h1c75;
aud[35648]=16'h1c62;
aud[35649]=16'h1c4e;
aud[35650]=16'h1c3b;
aud[35651]=16'h1c28;
aud[35652]=16'h1c15;
aud[35653]=16'h1c01;
aud[35654]=16'h1bee;
aud[35655]=16'h1bdb;
aud[35656]=16'h1bc8;
aud[35657]=16'h1bb4;
aud[35658]=16'h1ba1;
aud[35659]=16'h1b8d;
aud[35660]=16'h1b7a;
aud[35661]=16'h1b67;
aud[35662]=16'h1b53;
aud[35663]=16'h1b40;
aud[35664]=16'h1b2d;
aud[35665]=16'h1b19;
aud[35666]=16'h1b06;
aud[35667]=16'h1af2;
aud[35668]=16'h1adf;
aud[35669]=16'h1acb;
aud[35670]=16'h1ab8;
aud[35671]=16'h1aa4;
aud[35672]=16'h1a91;
aud[35673]=16'h1a7d;
aud[35674]=16'h1a6a;
aud[35675]=16'h1a56;
aud[35676]=16'h1a43;
aud[35677]=16'h1a2f;
aud[35678]=16'h1a1c;
aud[35679]=16'h1a08;
aud[35680]=16'h19f4;
aud[35681]=16'h19e1;
aud[35682]=16'h19cd;
aud[35683]=16'h19ba;
aud[35684]=16'h19a6;
aud[35685]=16'h1992;
aud[35686]=16'h197f;
aud[35687]=16'h196b;
aud[35688]=16'h1957;
aud[35689]=16'h1943;
aud[35690]=16'h1930;
aud[35691]=16'h191c;
aud[35692]=16'h1908;
aud[35693]=16'h18f5;
aud[35694]=16'h18e1;
aud[35695]=16'h18cd;
aud[35696]=16'h18b9;
aud[35697]=16'h18a5;
aud[35698]=16'h1892;
aud[35699]=16'h187e;
aud[35700]=16'h186a;
aud[35701]=16'h1856;
aud[35702]=16'h1842;
aud[35703]=16'h182f;
aud[35704]=16'h181b;
aud[35705]=16'h1807;
aud[35706]=16'h17f3;
aud[35707]=16'h17df;
aud[35708]=16'h17cb;
aud[35709]=16'h17b7;
aud[35710]=16'h17a3;
aud[35711]=16'h178f;
aud[35712]=16'h177b;
aud[35713]=16'h1767;
aud[35714]=16'h1753;
aud[35715]=16'h1740;
aud[35716]=16'h172c;
aud[35717]=16'h1718;
aud[35718]=16'h1704;
aud[35719]=16'h16f0;
aud[35720]=16'h16db;
aud[35721]=16'h16c7;
aud[35722]=16'h16b3;
aud[35723]=16'h169f;
aud[35724]=16'h168b;
aud[35725]=16'h1677;
aud[35726]=16'h1663;
aud[35727]=16'h164f;
aud[35728]=16'h163b;
aud[35729]=16'h1627;
aud[35730]=16'h1613;
aud[35731]=16'h15ff;
aud[35732]=16'h15ea;
aud[35733]=16'h15d6;
aud[35734]=16'h15c2;
aud[35735]=16'h15ae;
aud[35736]=16'h159a;
aud[35737]=16'h1586;
aud[35738]=16'h1571;
aud[35739]=16'h155d;
aud[35740]=16'h1549;
aud[35741]=16'h1535;
aud[35742]=16'h1520;
aud[35743]=16'h150c;
aud[35744]=16'h14f8;
aud[35745]=16'h14e4;
aud[35746]=16'h14cf;
aud[35747]=16'h14bb;
aud[35748]=16'h14a7;
aud[35749]=16'h1492;
aud[35750]=16'h147e;
aud[35751]=16'h146a;
aud[35752]=16'h1455;
aud[35753]=16'h1441;
aud[35754]=16'h142d;
aud[35755]=16'h1418;
aud[35756]=16'h1404;
aud[35757]=16'h13f0;
aud[35758]=16'h13db;
aud[35759]=16'h13c7;
aud[35760]=16'h13b3;
aud[35761]=16'h139e;
aud[35762]=16'h138a;
aud[35763]=16'h1375;
aud[35764]=16'h1361;
aud[35765]=16'h134c;
aud[35766]=16'h1338;
aud[35767]=16'h1323;
aud[35768]=16'h130f;
aud[35769]=16'h12fb;
aud[35770]=16'h12e6;
aud[35771]=16'h12d2;
aud[35772]=16'h12bd;
aud[35773]=16'h12a9;
aud[35774]=16'h1294;
aud[35775]=16'h127f;
aud[35776]=16'h126b;
aud[35777]=16'h1256;
aud[35778]=16'h1242;
aud[35779]=16'h122d;
aud[35780]=16'h1219;
aud[35781]=16'h1204;
aud[35782]=16'h11f0;
aud[35783]=16'h11db;
aud[35784]=16'h11c6;
aud[35785]=16'h11b2;
aud[35786]=16'h119d;
aud[35787]=16'h1189;
aud[35788]=16'h1174;
aud[35789]=16'h115f;
aud[35790]=16'h114b;
aud[35791]=16'h1136;
aud[35792]=16'h1121;
aud[35793]=16'h110d;
aud[35794]=16'h10f8;
aud[35795]=16'h10e3;
aud[35796]=16'h10cf;
aud[35797]=16'h10ba;
aud[35798]=16'h10a5;
aud[35799]=16'h1090;
aud[35800]=16'h107c;
aud[35801]=16'h1067;
aud[35802]=16'h1052;
aud[35803]=16'h103e;
aud[35804]=16'h1029;
aud[35805]=16'h1014;
aud[35806]=16'hfff;
aud[35807]=16'hfeb;
aud[35808]=16'hfd6;
aud[35809]=16'hfc1;
aud[35810]=16'hfac;
aud[35811]=16'hf97;
aud[35812]=16'hf83;
aud[35813]=16'hf6e;
aud[35814]=16'hf59;
aud[35815]=16'hf44;
aud[35816]=16'hf2f;
aud[35817]=16'hf1a;
aud[35818]=16'hf06;
aud[35819]=16'hef1;
aud[35820]=16'hedc;
aud[35821]=16'hec7;
aud[35822]=16'heb2;
aud[35823]=16'he9d;
aud[35824]=16'he88;
aud[35825]=16'he74;
aud[35826]=16'he5f;
aud[35827]=16'he4a;
aud[35828]=16'he35;
aud[35829]=16'he20;
aud[35830]=16'he0b;
aud[35831]=16'hdf6;
aud[35832]=16'hde1;
aud[35833]=16'hdcc;
aud[35834]=16'hdb7;
aud[35835]=16'hda2;
aud[35836]=16'hd8d;
aud[35837]=16'hd78;
aud[35838]=16'hd63;
aud[35839]=16'hd4e;
aud[35840]=16'hd39;
aud[35841]=16'hd24;
aud[35842]=16'hd0f;
aud[35843]=16'hcfa;
aud[35844]=16'hce5;
aud[35845]=16'hcd0;
aud[35846]=16'hcbb;
aud[35847]=16'hca6;
aud[35848]=16'hc91;
aud[35849]=16'hc7c;
aud[35850]=16'hc67;
aud[35851]=16'hc52;
aud[35852]=16'hc3d;
aud[35853]=16'hc28;
aud[35854]=16'hc13;
aud[35855]=16'hbfe;
aud[35856]=16'hbe9;
aud[35857]=16'hbd4;
aud[35858]=16'hbbf;
aud[35859]=16'hbaa;
aud[35860]=16'hb95;
aud[35861]=16'hb80;
aud[35862]=16'hb6a;
aud[35863]=16'hb55;
aud[35864]=16'hb40;
aud[35865]=16'hb2b;
aud[35866]=16'hb16;
aud[35867]=16'hb01;
aud[35868]=16'haec;
aud[35869]=16'had7;
aud[35870]=16'hac1;
aud[35871]=16'haac;
aud[35872]=16'ha97;
aud[35873]=16'ha82;
aud[35874]=16'ha6d;
aud[35875]=16'ha58;
aud[35876]=16'ha43;
aud[35877]=16'ha2d;
aud[35878]=16'ha18;
aud[35879]=16'ha03;
aud[35880]=16'h9ee;
aud[35881]=16'h9d9;
aud[35882]=16'h9c3;
aud[35883]=16'h9ae;
aud[35884]=16'h999;
aud[35885]=16'h984;
aud[35886]=16'h96f;
aud[35887]=16'h959;
aud[35888]=16'h944;
aud[35889]=16'h92f;
aud[35890]=16'h91a;
aud[35891]=16'h905;
aud[35892]=16'h8ef;
aud[35893]=16'h8da;
aud[35894]=16'h8c5;
aud[35895]=16'h8b0;
aud[35896]=16'h89a;
aud[35897]=16'h885;
aud[35898]=16'h870;
aud[35899]=16'h85b;
aud[35900]=16'h845;
aud[35901]=16'h830;
aud[35902]=16'h81b;
aud[35903]=16'h805;
aud[35904]=16'h7f0;
aud[35905]=16'h7db;
aud[35906]=16'h7c6;
aud[35907]=16'h7b0;
aud[35908]=16'h79b;
aud[35909]=16'h786;
aud[35910]=16'h770;
aud[35911]=16'h75b;
aud[35912]=16'h746;
aud[35913]=16'h731;
aud[35914]=16'h71b;
aud[35915]=16'h706;
aud[35916]=16'h6f1;
aud[35917]=16'h6db;
aud[35918]=16'h6c6;
aud[35919]=16'h6b1;
aud[35920]=16'h69b;
aud[35921]=16'h686;
aud[35922]=16'h671;
aud[35923]=16'h65b;
aud[35924]=16'h646;
aud[35925]=16'h631;
aud[35926]=16'h61b;
aud[35927]=16'h606;
aud[35928]=16'h5f1;
aud[35929]=16'h5db;
aud[35930]=16'h5c6;
aud[35931]=16'h5b0;
aud[35932]=16'h59b;
aud[35933]=16'h586;
aud[35934]=16'h570;
aud[35935]=16'h55b;
aud[35936]=16'h546;
aud[35937]=16'h530;
aud[35938]=16'h51b;
aud[35939]=16'h505;
aud[35940]=16'h4f0;
aud[35941]=16'h4db;
aud[35942]=16'h4c5;
aud[35943]=16'h4b0;
aud[35944]=16'h49b;
aud[35945]=16'h485;
aud[35946]=16'h470;
aud[35947]=16'h45a;
aud[35948]=16'h445;
aud[35949]=16'h430;
aud[35950]=16'h41a;
aud[35951]=16'h405;
aud[35952]=16'h3ef;
aud[35953]=16'h3da;
aud[35954]=16'h3c5;
aud[35955]=16'h3af;
aud[35956]=16'h39a;
aud[35957]=16'h384;
aud[35958]=16'h36f;
aud[35959]=16'h359;
aud[35960]=16'h344;
aud[35961]=16'h32f;
aud[35962]=16'h319;
aud[35963]=16'h304;
aud[35964]=16'h2ee;
aud[35965]=16'h2d9;
aud[35966]=16'h2c4;
aud[35967]=16'h2ae;
aud[35968]=16'h299;
aud[35969]=16'h283;
aud[35970]=16'h26e;
aud[35971]=16'h258;
aud[35972]=16'h243;
aud[35973]=16'h22e;
aud[35974]=16'h218;
aud[35975]=16'h203;
aud[35976]=16'h1ed;
aud[35977]=16'h1d8;
aud[35978]=16'h1c2;
aud[35979]=16'h1ad;
aud[35980]=16'h197;
aud[35981]=16'h182;
aud[35982]=16'h16d;
aud[35983]=16'h157;
aud[35984]=16'h142;
aud[35985]=16'h12c;
aud[35986]=16'h117;
aud[35987]=16'h101;
aud[35988]=16'hec;
aud[35989]=16'hd6;
aud[35990]=16'hc1;
aud[35991]=16'hac;
aud[35992]=16'h96;
aud[35993]=16'h81;
aud[35994]=16'h6b;
aud[35995]=16'h56;
aud[35996]=16'h40;
aud[35997]=16'h2b;
aud[35998]=16'h15;
aud[35999]=16'h0;
aud[36000]=16'hffeb;
aud[36001]=16'hffd5;
aud[36002]=16'hffc0;
aud[36003]=16'hffaa;
aud[36004]=16'hff95;
aud[36005]=16'hff7f;
aud[36006]=16'hff6a;
aud[36007]=16'hff54;
aud[36008]=16'hff3f;
aud[36009]=16'hff2a;
aud[36010]=16'hff14;
aud[36011]=16'hfeff;
aud[36012]=16'hfee9;
aud[36013]=16'hfed4;
aud[36014]=16'hfebe;
aud[36015]=16'hfea9;
aud[36016]=16'hfe93;
aud[36017]=16'hfe7e;
aud[36018]=16'hfe69;
aud[36019]=16'hfe53;
aud[36020]=16'hfe3e;
aud[36021]=16'hfe28;
aud[36022]=16'hfe13;
aud[36023]=16'hfdfd;
aud[36024]=16'hfde8;
aud[36025]=16'hfdd2;
aud[36026]=16'hfdbd;
aud[36027]=16'hfda8;
aud[36028]=16'hfd92;
aud[36029]=16'hfd7d;
aud[36030]=16'hfd67;
aud[36031]=16'hfd52;
aud[36032]=16'hfd3c;
aud[36033]=16'hfd27;
aud[36034]=16'hfd12;
aud[36035]=16'hfcfc;
aud[36036]=16'hfce7;
aud[36037]=16'hfcd1;
aud[36038]=16'hfcbc;
aud[36039]=16'hfca7;
aud[36040]=16'hfc91;
aud[36041]=16'hfc7c;
aud[36042]=16'hfc66;
aud[36043]=16'hfc51;
aud[36044]=16'hfc3b;
aud[36045]=16'hfc26;
aud[36046]=16'hfc11;
aud[36047]=16'hfbfb;
aud[36048]=16'hfbe6;
aud[36049]=16'hfbd0;
aud[36050]=16'hfbbb;
aud[36051]=16'hfba6;
aud[36052]=16'hfb90;
aud[36053]=16'hfb7b;
aud[36054]=16'hfb65;
aud[36055]=16'hfb50;
aud[36056]=16'hfb3b;
aud[36057]=16'hfb25;
aud[36058]=16'hfb10;
aud[36059]=16'hfafb;
aud[36060]=16'hfae5;
aud[36061]=16'hfad0;
aud[36062]=16'hfaba;
aud[36063]=16'hfaa5;
aud[36064]=16'hfa90;
aud[36065]=16'hfa7a;
aud[36066]=16'hfa65;
aud[36067]=16'hfa50;
aud[36068]=16'hfa3a;
aud[36069]=16'hfa25;
aud[36070]=16'hfa0f;
aud[36071]=16'hf9fa;
aud[36072]=16'hf9e5;
aud[36073]=16'hf9cf;
aud[36074]=16'hf9ba;
aud[36075]=16'hf9a5;
aud[36076]=16'hf98f;
aud[36077]=16'hf97a;
aud[36078]=16'hf965;
aud[36079]=16'hf94f;
aud[36080]=16'hf93a;
aud[36081]=16'hf925;
aud[36082]=16'hf90f;
aud[36083]=16'hf8fa;
aud[36084]=16'hf8e5;
aud[36085]=16'hf8cf;
aud[36086]=16'hf8ba;
aud[36087]=16'hf8a5;
aud[36088]=16'hf890;
aud[36089]=16'hf87a;
aud[36090]=16'hf865;
aud[36091]=16'hf850;
aud[36092]=16'hf83a;
aud[36093]=16'hf825;
aud[36094]=16'hf810;
aud[36095]=16'hf7fb;
aud[36096]=16'hf7e5;
aud[36097]=16'hf7d0;
aud[36098]=16'hf7bb;
aud[36099]=16'hf7a5;
aud[36100]=16'hf790;
aud[36101]=16'hf77b;
aud[36102]=16'hf766;
aud[36103]=16'hf750;
aud[36104]=16'hf73b;
aud[36105]=16'hf726;
aud[36106]=16'hf711;
aud[36107]=16'hf6fb;
aud[36108]=16'hf6e6;
aud[36109]=16'hf6d1;
aud[36110]=16'hf6bc;
aud[36111]=16'hf6a7;
aud[36112]=16'hf691;
aud[36113]=16'hf67c;
aud[36114]=16'hf667;
aud[36115]=16'hf652;
aud[36116]=16'hf63d;
aud[36117]=16'hf627;
aud[36118]=16'hf612;
aud[36119]=16'hf5fd;
aud[36120]=16'hf5e8;
aud[36121]=16'hf5d3;
aud[36122]=16'hf5bd;
aud[36123]=16'hf5a8;
aud[36124]=16'hf593;
aud[36125]=16'hf57e;
aud[36126]=16'hf569;
aud[36127]=16'hf554;
aud[36128]=16'hf53f;
aud[36129]=16'hf529;
aud[36130]=16'hf514;
aud[36131]=16'hf4ff;
aud[36132]=16'hf4ea;
aud[36133]=16'hf4d5;
aud[36134]=16'hf4c0;
aud[36135]=16'hf4ab;
aud[36136]=16'hf496;
aud[36137]=16'hf480;
aud[36138]=16'hf46b;
aud[36139]=16'hf456;
aud[36140]=16'hf441;
aud[36141]=16'hf42c;
aud[36142]=16'hf417;
aud[36143]=16'hf402;
aud[36144]=16'hf3ed;
aud[36145]=16'hf3d8;
aud[36146]=16'hf3c3;
aud[36147]=16'hf3ae;
aud[36148]=16'hf399;
aud[36149]=16'hf384;
aud[36150]=16'hf36f;
aud[36151]=16'hf35a;
aud[36152]=16'hf345;
aud[36153]=16'hf330;
aud[36154]=16'hf31b;
aud[36155]=16'hf306;
aud[36156]=16'hf2f1;
aud[36157]=16'hf2dc;
aud[36158]=16'hf2c7;
aud[36159]=16'hf2b2;
aud[36160]=16'hf29d;
aud[36161]=16'hf288;
aud[36162]=16'hf273;
aud[36163]=16'hf25e;
aud[36164]=16'hf249;
aud[36165]=16'hf234;
aud[36166]=16'hf21f;
aud[36167]=16'hf20a;
aud[36168]=16'hf1f5;
aud[36169]=16'hf1e0;
aud[36170]=16'hf1cb;
aud[36171]=16'hf1b6;
aud[36172]=16'hf1a1;
aud[36173]=16'hf18c;
aud[36174]=16'hf178;
aud[36175]=16'hf163;
aud[36176]=16'hf14e;
aud[36177]=16'hf139;
aud[36178]=16'hf124;
aud[36179]=16'hf10f;
aud[36180]=16'hf0fa;
aud[36181]=16'hf0e6;
aud[36182]=16'hf0d1;
aud[36183]=16'hf0bc;
aud[36184]=16'hf0a7;
aud[36185]=16'hf092;
aud[36186]=16'hf07d;
aud[36187]=16'hf069;
aud[36188]=16'hf054;
aud[36189]=16'hf03f;
aud[36190]=16'hf02a;
aud[36191]=16'hf015;
aud[36192]=16'hf001;
aud[36193]=16'hefec;
aud[36194]=16'hefd7;
aud[36195]=16'hefc2;
aud[36196]=16'hefae;
aud[36197]=16'hef99;
aud[36198]=16'hef84;
aud[36199]=16'hef70;
aud[36200]=16'hef5b;
aud[36201]=16'hef46;
aud[36202]=16'hef31;
aud[36203]=16'hef1d;
aud[36204]=16'hef08;
aud[36205]=16'heef3;
aud[36206]=16'heedf;
aud[36207]=16'heeca;
aud[36208]=16'heeb5;
aud[36209]=16'heea1;
aud[36210]=16'hee8c;
aud[36211]=16'hee77;
aud[36212]=16'hee63;
aud[36213]=16'hee4e;
aud[36214]=16'hee3a;
aud[36215]=16'hee25;
aud[36216]=16'hee10;
aud[36217]=16'hedfc;
aud[36218]=16'hede7;
aud[36219]=16'hedd3;
aud[36220]=16'hedbe;
aud[36221]=16'hedaa;
aud[36222]=16'hed95;
aud[36223]=16'hed81;
aud[36224]=16'hed6c;
aud[36225]=16'hed57;
aud[36226]=16'hed43;
aud[36227]=16'hed2e;
aud[36228]=16'hed1a;
aud[36229]=16'hed05;
aud[36230]=16'hecf1;
aud[36231]=16'hecdd;
aud[36232]=16'hecc8;
aud[36233]=16'hecb4;
aud[36234]=16'hec9f;
aud[36235]=16'hec8b;
aud[36236]=16'hec76;
aud[36237]=16'hec62;
aud[36238]=16'hec4d;
aud[36239]=16'hec39;
aud[36240]=16'hec25;
aud[36241]=16'hec10;
aud[36242]=16'hebfc;
aud[36243]=16'hebe8;
aud[36244]=16'hebd3;
aud[36245]=16'hebbf;
aud[36246]=16'hebab;
aud[36247]=16'heb96;
aud[36248]=16'heb82;
aud[36249]=16'heb6e;
aud[36250]=16'heb59;
aud[36251]=16'heb45;
aud[36252]=16'heb31;
aud[36253]=16'heb1c;
aud[36254]=16'heb08;
aud[36255]=16'heaf4;
aud[36256]=16'heae0;
aud[36257]=16'heacb;
aud[36258]=16'heab7;
aud[36259]=16'heaa3;
aud[36260]=16'hea8f;
aud[36261]=16'hea7a;
aud[36262]=16'hea66;
aud[36263]=16'hea52;
aud[36264]=16'hea3e;
aud[36265]=16'hea2a;
aud[36266]=16'hea16;
aud[36267]=16'hea01;
aud[36268]=16'he9ed;
aud[36269]=16'he9d9;
aud[36270]=16'he9c5;
aud[36271]=16'he9b1;
aud[36272]=16'he99d;
aud[36273]=16'he989;
aud[36274]=16'he975;
aud[36275]=16'he961;
aud[36276]=16'he94d;
aud[36277]=16'he939;
aud[36278]=16'he925;
aud[36279]=16'he910;
aud[36280]=16'he8fc;
aud[36281]=16'he8e8;
aud[36282]=16'he8d4;
aud[36283]=16'he8c0;
aud[36284]=16'he8ad;
aud[36285]=16'he899;
aud[36286]=16'he885;
aud[36287]=16'he871;
aud[36288]=16'he85d;
aud[36289]=16'he849;
aud[36290]=16'he835;
aud[36291]=16'he821;
aud[36292]=16'he80d;
aud[36293]=16'he7f9;
aud[36294]=16'he7e5;
aud[36295]=16'he7d1;
aud[36296]=16'he7be;
aud[36297]=16'he7aa;
aud[36298]=16'he796;
aud[36299]=16'he782;
aud[36300]=16'he76e;
aud[36301]=16'he75b;
aud[36302]=16'he747;
aud[36303]=16'he733;
aud[36304]=16'he71f;
aud[36305]=16'he70b;
aud[36306]=16'he6f8;
aud[36307]=16'he6e4;
aud[36308]=16'he6d0;
aud[36309]=16'he6bd;
aud[36310]=16'he6a9;
aud[36311]=16'he695;
aud[36312]=16'he681;
aud[36313]=16'he66e;
aud[36314]=16'he65a;
aud[36315]=16'he646;
aud[36316]=16'he633;
aud[36317]=16'he61f;
aud[36318]=16'he60c;
aud[36319]=16'he5f8;
aud[36320]=16'he5e4;
aud[36321]=16'he5d1;
aud[36322]=16'he5bd;
aud[36323]=16'he5aa;
aud[36324]=16'he596;
aud[36325]=16'he583;
aud[36326]=16'he56f;
aud[36327]=16'he55c;
aud[36328]=16'he548;
aud[36329]=16'he535;
aud[36330]=16'he521;
aud[36331]=16'he50e;
aud[36332]=16'he4fa;
aud[36333]=16'he4e7;
aud[36334]=16'he4d3;
aud[36335]=16'he4c0;
aud[36336]=16'he4ad;
aud[36337]=16'he499;
aud[36338]=16'he486;
aud[36339]=16'he473;
aud[36340]=16'he45f;
aud[36341]=16'he44c;
aud[36342]=16'he438;
aud[36343]=16'he425;
aud[36344]=16'he412;
aud[36345]=16'he3ff;
aud[36346]=16'he3eb;
aud[36347]=16'he3d8;
aud[36348]=16'he3c5;
aud[36349]=16'he3b2;
aud[36350]=16'he39e;
aud[36351]=16'he38b;
aud[36352]=16'he378;
aud[36353]=16'he365;
aud[36354]=16'he352;
aud[36355]=16'he33e;
aud[36356]=16'he32b;
aud[36357]=16'he318;
aud[36358]=16'he305;
aud[36359]=16'he2f2;
aud[36360]=16'he2df;
aud[36361]=16'he2cc;
aud[36362]=16'he2b9;
aud[36363]=16'he2a5;
aud[36364]=16'he292;
aud[36365]=16'he27f;
aud[36366]=16'he26c;
aud[36367]=16'he259;
aud[36368]=16'he246;
aud[36369]=16'he233;
aud[36370]=16'he220;
aud[36371]=16'he20d;
aud[36372]=16'he1fa;
aud[36373]=16'he1e8;
aud[36374]=16'he1d5;
aud[36375]=16'he1c2;
aud[36376]=16'he1af;
aud[36377]=16'he19c;
aud[36378]=16'he189;
aud[36379]=16'he176;
aud[36380]=16'he163;
aud[36381]=16'he151;
aud[36382]=16'he13e;
aud[36383]=16'he12b;
aud[36384]=16'he118;
aud[36385]=16'he105;
aud[36386]=16'he0f3;
aud[36387]=16'he0e0;
aud[36388]=16'he0cd;
aud[36389]=16'he0ba;
aud[36390]=16'he0a8;
aud[36391]=16'he095;
aud[36392]=16'he082;
aud[36393]=16'he070;
aud[36394]=16'he05d;
aud[36395]=16'he04a;
aud[36396]=16'he038;
aud[36397]=16'he025;
aud[36398]=16'he013;
aud[36399]=16'he000;
aud[36400]=16'hdfed;
aud[36401]=16'hdfdb;
aud[36402]=16'hdfc8;
aud[36403]=16'hdfb6;
aud[36404]=16'hdfa3;
aud[36405]=16'hdf91;
aud[36406]=16'hdf7e;
aud[36407]=16'hdf6c;
aud[36408]=16'hdf59;
aud[36409]=16'hdf47;
aud[36410]=16'hdf35;
aud[36411]=16'hdf22;
aud[36412]=16'hdf10;
aud[36413]=16'hdefd;
aud[36414]=16'hdeeb;
aud[36415]=16'hded9;
aud[36416]=16'hdec6;
aud[36417]=16'hdeb4;
aud[36418]=16'hdea2;
aud[36419]=16'hde8f;
aud[36420]=16'hde7d;
aud[36421]=16'hde6b;
aud[36422]=16'hde59;
aud[36423]=16'hde46;
aud[36424]=16'hde34;
aud[36425]=16'hde22;
aud[36426]=16'hde10;
aud[36427]=16'hddfe;
aud[36428]=16'hddeb;
aud[36429]=16'hddd9;
aud[36430]=16'hddc7;
aud[36431]=16'hddb5;
aud[36432]=16'hdda3;
aud[36433]=16'hdd91;
aud[36434]=16'hdd7f;
aud[36435]=16'hdd6d;
aud[36436]=16'hdd5b;
aud[36437]=16'hdd49;
aud[36438]=16'hdd37;
aud[36439]=16'hdd25;
aud[36440]=16'hdd13;
aud[36441]=16'hdd01;
aud[36442]=16'hdcef;
aud[36443]=16'hdcdd;
aud[36444]=16'hdccb;
aud[36445]=16'hdcb9;
aud[36446]=16'hdca7;
aud[36447]=16'hdc95;
aud[36448]=16'hdc83;
aud[36449]=16'hdc72;
aud[36450]=16'hdc60;
aud[36451]=16'hdc4e;
aud[36452]=16'hdc3c;
aud[36453]=16'hdc2a;
aud[36454]=16'hdc19;
aud[36455]=16'hdc07;
aud[36456]=16'hdbf5;
aud[36457]=16'hdbe3;
aud[36458]=16'hdbd2;
aud[36459]=16'hdbc0;
aud[36460]=16'hdbae;
aud[36461]=16'hdb9d;
aud[36462]=16'hdb8b;
aud[36463]=16'hdb79;
aud[36464]=16'hdb68;
aud[36465]=16'hdb56;
aud[36466]=16'hdb45;
aud[36467]=16'hdb33;
aud[36468]=16'hdb22;
aud[36469]=16'hdb10;
aud[36470]=16'hdaff;
aud[36471]=16'hdaed;
aud[36472]=16'hdadc;
aud[36473]=16'hdaca;
aud[36474]=16'hdab9;
aud[36475]=16'hdaa7;
aud[36476]=16'hda96;
aud[36477]=16'hda84;
aud[36478]=16'hda73;
aud[36479]=16'hda62;
aud[36480]=16'hda50;
aud[36481]=16'hda3f;
aud[36482]=16'hda2e;
aud[36483]=16'hda1c;
aud[36484]=16'hda0b;
aud[36485]=16'hd9fa;
aud[36486]=16'hd9e9;
aud[36487]=16'hd9d7;
aud[36488]=16'hd9c6;
aud[36489]=16'hd9b5;
aud[36490]=16'hd9a4;
aud[36491]=16'hd993;
aud[36492]=16'hd982;
aud[36493]=16'hd970;
aud[36494]=16'hd95f;
aud[36495]=16'hd94e;
aud[36496]=16'hd93d;
aud[36497]=16'hd92c;
aud[36498]=16'hd91b;
aud[36499]=16'hd90a;
aud[36500]=16'hd8f9;
aud[36501]=16'hd8e8;
aud[36502]=16'hd8d7;
aud[36503]=16'hd8c6;
aud[36504]=16'hd8b5;
aud[36505]=16'hd8a4;
aud[36506]=16'hd893;
aud[36507]=16'hd882;
aud[36508]=16'hd872;
aud[36509]=16'hd861;
aud[36510]=16'hd850;
aud[36511]=16'hd83f;
aud[36512]=16'hd82e;
aud[36513]=16'hd81e;
aud[36514]=16'hd80d;
aud[36515]=16'hd7fc;
aud[36516]=16'hd7eb;
aud[36517]=16'hd7db;
aud[36518]=16'hd7ca;
aud[36519]=16'hd7b9;
aud[36520]=16'hd7a9;
aud[36521]=16'hd798;
aud[36522]=16'hd787;
aud[36523]=16'hd777;
aud[36524]=16'hd766;
aud[36525]=16'hd756;
aud[36526]=16'hd745;
aud[36527]=16'hd734;
aud[36528]=16'hd724;
aud[36529]=16'hd713;
aud[36530]=16'hd703;
aud[36531]=16'hd6f2;
aud[36532]=16'hd6e2;
aud[36533]=16'hd6d2;
aud[36534]=16'hd6c1;
aud[36535]=16'hd6b1;
aud[36536]=16'hd6a0;
aud[36537]=16'hd690;
aud[36538]=16'hd680;
aud[36539]=16'hd66f;
aud[36540]=16'hd65f;
aud[36541]=16'hd64f;
aud[36542]=16'hd63f;
aud[36543]=16'hd62e;
aud[36544]=16'hd61e;
aud[36545]=16'hd60e;
aud[36546]=16'hd5fe;
aud[36547]=16'hd5ee;
aud[36548]=16'hd5dd;
aud[36549]=16'hd5cd;
aud[36550]=16'hd5bd;
aud[36551]=16'hd5ad;
aud[36552]=16'hd59d;
aud[36553]=16'hd58d;
aud[36554]=16'hd57d;
aud[36555]=16'hd56d;
aud[36556]=16'hd55d;
aud[36557]=16'hd54d;
aud[36558]=16'hd53d;
aud[36559]=16'hd52d;
aud[36560]=16'hd51d;
aud[36561]=16'hd50d;
aud[36562]=16'hd4fd;
aud[36563]=16'hd4ed;
aud[36564]=16'hd4de;
aud[36565]=16'hd4ce;
aud[36566]=16'hd4be;
aud[36567]=16'hd4ae;
aud[36568]=16'hd49e;
aud[36569]=16'hd48f;
aud[36570]=16'hd47f;
aud[36571]=16'hd46f;
aud[36572]=16'hd45f;
aud[36573]=16'hd450;
aud[36574]=16'hd440;
aud[36575]=16'hd430;
aud[36576]=16'hd421;
aud[36577]=16'hd411;
aud[36578]=16'hd402;
aud[36579]=16'hd3f2;
aud[36580]=16'hd3e2;
aud[36581]=16'hd3d3;
aud[36582]=16'hd3c3;
aud[36583]=16'hd3b4;
aud[36584]=16'hd3a4;
aud[36585]=16'hd395;
aud[36586]=16'hd386;
aud[36587]=16'hd376;
aud[36588]=16'hd367;
aud[36589]=16'hd357;
aud[36590]=16'hd348;
aud[36591]=16'hd339;
aud[36592]=16'hd329;
aud[36593]=16'hd31a;
aud[36594]=16'hd30b;
aud[36595]=16'hd2fc;
aud[36596]=16'hd2ec;
aud[36597]=16'hd2dd;
aud[36598]=16'hd2ce;
aud[36599]=16'hd2bf;
aud[36600]=16'hd2b0;
aud[36601]=16'hd2a0;
aud[36602]=16'hd291;
aud[36603]=16'hd282;
aud[36604]=16'hd273;
aud[36605]=16'hd264;
aud[36606]=16'hd255;
aud[36607]=16'hd246;
aud[36608]=16'hd237;
aud[36609]=16'hd228;
aud[36610]=16'hd219;
aud[36611]=16'hd20a;
aud[36612]=16'hd1fb;
aud[36613]=16'hd1ec;
aud[36614]=16'hd1de;
aud[36615]=16'hd1cf;
aud[36616]=16'hd1c0;
aud[36617]=16'hd1b1;
aud[36618]=16'hd1a2;
aud[36619]=16'hd193;
aud[36620]=16'hd185;
aud[36621]=16'hd176;
aud[36622]=16'hd167;
aud[36623]=16'hd159;
aud[36624]=16'hd14a;
aud[36625]=16'hd13b;
aud[36626]=16'hd12d;
aud[36627]=16'hd11e;
aud[36628]=16'hd10f;
aud[36629]=16'hd101;
aud[36630]=16'hd0f2;
aud[36631]=16'hd0e4;
aud[36632]=16'hd0d5;
aud[36633]=16'hd0c7;
aud[36634]=16'hd0b8;
aud[36635]=16'hd0aa;
aud[36636]=16'hd09b;
aud[36637]=16'hd08d;
aud[36638]=16'hd07f;
aud[36639]=16'hd070;
aud[36640]=16'hd062;
aud[36641]=16'hd054;
aud[36642]=16'hd045;
aud[36643]=16'hd037;
aud[36644]=16'hd029;
aud[36645]=16'hd01b;
aud[36646]=16'hd00c;
aud[36647]=16'hcffe;
aud[36648]=16'hcff0;
aud[36649]=16'hcfe2;
aud[36650]=16'hcfd4;
aud[36651]=16'hcfc6;
aud[36652]=16'hcfb8;
aud[36653]=16'hcfa9;
aud[36654]=16'hcf9b;
aud[36655]=16'hcf8d;
aud[36656]=16'hcf7f;
aud[36657]=16'hcf71;
aud[36658]=16'hcf63;
aud[36659]=16'hcf56;
aud[36660]=16'hcf48;
aud[36661]=16'hcf3a;
aud[36662]=16'hcf2c;
aud[36663]=16'hcf1e;
aud[36664]=16'hcf10;
aud[36665]=16'hcf02;
aud[36666]=16'hcef5;
aud[36667]=16'hcee7;
aud[36668]=16'hced9;
aud[36669]=16'hcecb;
aud[36670]=16'hcebe;
aud[36671]=16'hceb0;
aud[36672]=16'hcea2;
aud[36673]=16'hce95;
aud[36674]=16'hce87;
aud[36675]=16'hce79;
aud[36676]=16'hce6c;
aud[36677]=16'hce5e;
aud[36678]=16'hce51;
aud[36679]=16'hce43;
aud[36680]=16'hce36;
aud[36681]=16'hce28;
aud[36682]=16'hce1b;
aud[36683]=16'hce0d;
aud[36684]=16'hce00;
aud[36685]=16'hcdf3;
aud[36686]=16'hcde5;
aud[36687]=16'hcdd8;
aud[36688]=16'hcdcb;
aud[36689]=16'hcdbd;
aud[36690]=16'hcdb0;
aud[36691]=16'hcda3;
aud[36692]=16'hcd96;
aud[36693]=16'hcd88;
aud[36694]=16'hcd7b;
aud[36695]=16'hcd6e;
aud[36696]=16'hcd61;
aud[36697]=16'hcd54;
aud[36698]=16'hcd47;
aud[36699]=16'hcd3a;
aud[36700]=16'hcd2d;
aud[36701]=16'hcd20;
aud[36702]=16'hcd13;
aud[36703]=16'hcd06;
aud[36704]=16'hccf9;
aud[36705]=16'hccec;
aud[36706]=16'hccdf;
aud[36707]=16'hccd2;
aud[36708]=16'hccc5;
aud[36709]=16'hccb8;
aud[36710]=16'hccab;
aud[36711]=16'hcc9f;
aud[36712]=16'hcc92;
aud[36713]=16'hcc85;
aud[36714]=16'hcc78;
aud[36715]=16'hcc6c;
aud[36716]=16'hcc5f;
aud[36717]=16'hcc52;
aud[36718]=16'hcc46;
aud[36719]=16'hcc39;
aud[36720]=16'hcc2c;
aud[36721]=16'hcc20;
aud[36722]=16'hcc13;
aud[36723]=16'hcc07;
aud[36724]=16'hcbfa;
aud[36725]=16'hcbee;
aud[36726]=16'hcbe1;
aud[36727]=16'hcbd5;
aud[36728]=16'hcbc9;
aud[36729]=16'hcbbc;
aud[36730]=16'hcbb0;
aud[36731]=16'hcba3;
aud[36732]=16'hcb97;
aud[36733]=16'hcb8b;
aud[36734]=16'hcb7f;
aud[36735]=16'hcb72;
aud[36736]=16'hcb66;
aud[36737]=16'hcb5a;
aud[36738]=16'hcb4e;
aud[36739]=16'hcb42;
aud[36740]=16'hcb35;
aud[36741]=16'hcb29;
aud[36742]=16'hcb1d;
aud[36743]=16'hcb11;
aud[36744]=16'hcb05;
aud[36745]=16'hcaf9;
aud[36746]=16'hcaed;
aud[36747]=16'hcae1;
aud[36748]=16'hcad5;
aud[36749]=16'hcac9;
aud[36750]=16'hcabd;
aud[36751]=16'hcab1;
aud[36752]=16'hcaa6;
aud[36753]=16'hca9a;
aud[36754]=16'hca8e;
aud[36755]=16'hca82;
aud[36756]=16'hca76;
aud[36757]=16'hca6b;
aud[36758]=16'hca5f;
aud[36759]=16'hca53;
aud[36760]=16'hca48;
aud[36761]=16'hca3c;
aud[36762]=16'hca30;
aud[36763]=16'hca25;
aud[36764]=16'hca19;
aud[36765]=16'hca0e;
aud[36766]=16'hca02;
aud[36767]=16'hc9f7;
aud[36768]=16'hc9eb;
aud[36769]=16'hc9e0;
aud[36770]=16'hc9d4;
aud[36771]=16'hc9c9;
aud[36772]=16'hc9bd;
aud[36773]=16'hc9b2;
aud[36774]=16'hc9a7;
aud[36775]=16'hc99b;
aud[36776]=16'hc990;
aud[36777]=16'hc985;
aud[36778]=16'hc97a;
aud[36779]=16'hc96e;
aud[36780]=16'hc963;
aud[36781]=16'hc958;
aud[36782]=16'hc94d;
aud[36783]=16'hc942;
aud[36784]=16'hc937;
aud[36785]=16'hc92c;
aud[36786]=16'hc920;
aud[36787]=16'hc915;
aud[36788]=16'hc90a;
aud[36789]=16'hc8ff;
aud[36790]=16'hc8f5;
aud[36791]=16'hc8ea;
aud[36792]=16'hc8df;
aud[36793]=16'hc8d4;
aud[36794]=16'hc8c9;
aud[36795]=16'hc8be;
aud[36796]=16'hc8b3;
aud[36797]=16'hc8a9;
aud[36798]=16'hc89e;
aud[36799]=16'hc893;
aud[36800]=16'hc888;
aud[36801]=16'hc87e;
aud[36802]=16'hc873;
aud[36803]=16'hc868;
aud[36804]=16'hc85e;
aud[36805]=16'hc853;
aud[36806]=16'hc849;
aud[36807]=16'hc83e;
aud[36808]=16'hc834;
aud[36809]=16'hc829;
aud[36810]=16'hc81f;
aud[36811]=16'hc814;
aud[36812]=16'hc80a;
aud[36813]=16'hc7ff;
aud[36814]=16'hc7f5;
aud[36815]=16'hc7eb;
aud[36816]=16'hc7e0;
aud[36817]=16'hc7d6;
aud[36818]=16'hc7cc;
aud[36819]=16'hc7c1;
aud[36820]=16'hc7b7;
aud[36821]=16'hc7ad;
aud[36822]=16'hc7a3;
aud[36823]=16'hc799;
aud[36824]=16'hc78f;
aud[36825]=16'hc785;
aud[36826]=16'hc77a;
aud[36827]=16'hc770;
aud[36828]=16'hc766;
aud[36829]=16'hc75c;
aud[36830]=16'hc752;
aud[36831]=16'hc748;
aud[36832]=16'hc73f;
aud[36833]=16'hc735;
aud[36834]=16'hc72b;
aud[36835]=16'hc721;
aud[36836]=16'hc717;
aud[36837]=16'hc70d;
aud[36838]=16'hc703;
aud[36839]=16'hc6fa;
aud[36840]=16'hc6f0;
aud[36841]=16'hc6e6;
aud[36842]=16'hc6dd;
aud[36843]=16'hc6d3;
aud[36844]=16'hc6c9;
aud[36845]=16'hc6c0;
aud[36846]=16'hc6b6;
aud[36847]=16'hc6ad;
aud[36848]=16'hc6a3;
aud[36849]=16'hc69a;
aud[36850]=16'hc690;
aud[36851]=16'hc687;
aud[36852]=16'hc67d;
aud[36853]=16'hc674;
aud[36854]=16'hc66b;
aud[36855]=16'hc661;
aud[36856]=16'hc658;
aud[36857]=16'hc64f;
aud[36858]=16'hc645;
aud[36859]=16'hc63c;
aud[36860]=16'hc633;
aud[36861]=16'hc62a;
aud[36862]=16'hc620;
aud[36863]=16'hc617;
aud[36864]=16'hc60e;
aud[36865]=16'hc605;
aud[36866]=16'hc5fc;
aud[36867]=16'hc5f3;
aud[36868]=16'hc5ea;
aud[36869]=16'hc5e1;
aud[36870]=16'hc5d8;
aud[36871]=16'hc5cf;
aud[36872]=16'hc5c6;
aud[36873]=16'hc5bd;
aud[36874]=16'hc5b4;
aud[36875]=16'hc5ac;
aud[36876]=16'hc5a3;
aud[36877]=16'hc59a;
aud[36878]=16'hc591;
aud[36879]=16'hc588;
aud[36880]=16'hc580;
aud[36881]=16'hc577;
aud[36882]=16'hc56e;
aud[36883]=16'hc566;
aud[36884]=16'hc55d;
aud[36885]=16'hc555;
aud[36886]=16'hc54c;
aud[36887]=16'hc544;
aud[36888]=16'hc53b;
aud[36889]=16'hc533;
aud[36890]=16'hc52a;
aud[36891]=16'hc522;
aud[36892]=16'hc519;
aud[36893]=16'hc511;
aud[36894]=16'hc509;
aud[36895]=16'hc500;
aud[36896]=16'hc4f8;
aud[36897]=16'hc4f0;
aud[36898]=16'hc4e7;
aud[36899]=16'hc4df;
aud[36900]=16'hc4d7;
aud[36901]=16'hc4cf;
aud[36902]=16'hc4c7;
aud[36903]=16'hc4bf;
aud[36904]=16'hc4b6;
aud[36905]=16'hc4ae;
aud[36906]=16'hc4a6;
aud[36907]=16'hc49e;
aud[36908]=16'hc496;
aud[36909]=16'hc48e;
aud[36910]=16'hc486;
aud[36911]=16'hc47f;
aud[36912]=16'hc477;
aud[36913]=16'hc46f;
aud[36914]=16'hc467;
aud[36915]=16'hc45f;
aud[36916]=16'hc457;
aud[36917]=16'hc450;
aud[36918]=16'hc448;
aud[36919]=16'hc440;
aud[36920]=16'hc439;
aud[36921]=16'hc431;
aud[36922]=16'hc429;
aud[36923]=16'hc422;
aud[36924]=16'hc41a;
aud[36925]=16'hc413;
aud[36926]=16'hc40b;
aud[36927]=16'hc404;
aud[36928]=16'hc3fc;
aud[36929]=16'hc3f5;
aud[36930]=16'hc3ed;
aud[36931]=16'hc3e6;
aud[36932]=16'hc3df;
aud[36933]=16'hc3d7;
aud[36934]=16'hc3d0;
aud[36935]=16'hc3c9;
aud[36936]=16'hc3c1;
aud[36937]=16'hc3ba;
aud[36938]=16'hc3b3;
aud[36939]=16'hc3ac;
aud[36940]=16'hc3a5;
aud[36941]=16'hc39d;
aud[36942]=16'hc396;
aud[36943]=16'hc38f;
aud[36944]=16'hc388;
aud[36945]=16'hc381;
aud[36946]=16'hc37a;
aud[36947]=16'hc373;
aud[36948]=16'hc36c;
aud[36949]=16'hc365;
aud[36950]=16'hc35f;
aud[36951]=16'hc358;
aud[36952]=16'hc351;
aud[36953]=16'hc34a;
aud[36954]=16'hc343;
aud[36955]=16'hc33d;
aud[36956]=16'hc336;
aud[36957]=16'hc32f;
aud[36958]=16'hc329;
aud[36959]=16'hc322;
aud[36960]=16'hc31b;
aud[36961]=16'hc315;
aud[36962]=16'hc30e;
aud[36963]=16'hc308;
aud[36964]=16'hc301;
aud[36965]=16'hc2fb;
aud[36966]=16'hc2f4;
aud[36967]=16'hc2ee;
aud[36968]=16'hc2e7;
aud[36969]=16'hc2e1;
aud[36970]=16'hc2db;
aud[36971]=16'hc2d4;
aud[36972]=16'hc2ce;
aud[36973]=16'hc2c8;
aud[36974]=16'hc2c1;
aud[36975]=16'hc2bb;
aud[36976]=16'hc2b5;
aud[36977]=16'hc2af;
aud[36978]=16'hc2a9;
aud[36979]=16'hc2a3;
aud[36980]=16'hc29d;
aud[36981]=16'hc297;
aud[36982]=16'hc291;
aud[36983]=16'hc28b;
aud[36984]=16'hc285;
aud[36985]=16'hc27f;
aud[36986]=16'hc279;
aud[36987]=16'hc273;
aud[36988]=16'hc26d;
aud[36989]=16'hc267;
aud[36990]=16'hc261;
aud[36991]=16'hc25c;
aud[36992]=16'hc256;
aud[36993]=16'hc250;
aud[36994]=16'hc24a;
aud[36995]=16'hc245;
aud[36996]=16'hc23f;
aud[36997]=16'hc239;
aud[36998]=16'hc234;
aud[36999]=16'hc22e;
aud[37000]=16'hc229;
aud[37001]=16'hc223;
aud[37002]=16'hc21e;
aud[37003]=16'hc218;
aud[37004]=16'hc213;
aud[37005]=16'hc20d;
aud[37006]=16'hc208;
aud[37007]=16'hc203;
aud[37008]=16'hc1fd;
aud[37009]=16'hc1f8;
aud[37010]=16'hc1f3;
aud[37011]=16'hc1ee;
aud[37012]=16'hc1e8;
aud[37013]=16'hc1e3;
aud[37014]=16'hc1de;
aud[37015]=16'hc1d9;
aud[37016]=16'hc1d4;
aud[37017]=16'hc1cf;
aud[37018]=16'hc1ca;
aud[37019]=16'hc1c5;
aud[37020]=16'hc1c0;
aud[37021]=16'hc1bb;
aud[37022]=16'hc1b6;
aud[37023]=16'hc1b1;
aud[37024]=16'hc1ac;
aud[37025]=16'hc1a7;
aud[37026]=16'hc1a2;
aud[37027]=16'hc19e;
aud[37028]=16'hc199;
aud[37029]=16'hc194;
aud[37030]=16'hc18f;
aud[37031]=16'hc18b;
aud[37032]=16'hc186;
aud[37033]=16'hc181;
aud[37034]=16'hc17d;
aud[37035]=16'hc178;
aud[37036]=16'hc174;
aud[37037]=16'hc16f;
aud[37038]=16'hc16b;
aud[37039]=16'hc166;
aud[37040]=16'hc162;
aud[37041]=16'hc15d;
aud[37042]=16'hc159;
aud[37043]=16'hc154;
aud[37044]=16'hc150;
aud[37045]=16'hc14c;
aud[37046]=16'hc147;
aud[37047]=16'hc143;
aud[37048]=16'hc13f;
aud[37049]=16'hc13b;
aud[37050]=16'hc137;
aud[37051]=16'hc133;
aud[37052]=16'hc12e;
aud[37053]=16'hc12a;
aud[37054]=16'hc126;
aud[37055]=16'hc122;
aud[37056]=16'hc11e;
aud[37057]=16'hc11a;
aud[37058]=16'hc116;
aud[37059]=16'hc112;
aud[37060]=16'hc10e;
aud[37061]=16'hc10b;
aud[37062]=16'hc107;
aud[37063]=16'hc103;
aud[37064]=16'hc0ff;
aud[37065]=16'hc0fb;
aud[37066]=16'hc0f8;
aud[37067]=16'hc0f4;
aud[37068]=16'hc0f0;
aud[37069]=16'hc0ed;
aud[37070]=16'hc0e9;
aud[37071]=16'hc0e5;
aud[37072]=16'hc0e2;
aud[37073]=16'hc0de;
aud[37074]=16'hc0db;
aud[37075]=16'hc0d7;
aud[37076]=16'hc0d4;
aud[37077]=16'hc0d0;
aud[37078]=16'hc0cd;
aud[37079]=16'hc0ca;
aud[37080]=16'hc0c6;
aud[37081]=16'hc0c3;
aud[37082]=16'hc0c0;
aud[37083]=16'hc0bd;
aud[37084]=16'hc0b9;
aud[37085]=16'hc0b6;
aud[37086]=16'hc0b3;
aud[37087]=16'hc0b0;
aud[37088]=16'hc0ad;
aud[37089]=16'hc0aa;
aud[37090]=16'hc0a6;
aud[37091]=16'hc0a3;
aud[37092]=16'hc0a0;
aud[37093]=16'hc09d;
aud[37094]=16'hc09b;
aud[37095]=16'hc098;
aud[37096]=16'hc095;
aud[37097]=16'hc092;
aud[37098]=16'hc08f;
aud[37099]=16'hc08c;
aud[37100]=16'hc089;
aud[37101]=16'hc087;
aud[37102]=16'hc084;
aud[37103]=16'hc081;
aud[37104]=16'hc07f;
aud[37105]=16'hc07c;
aud[37106]=16'hc079;
aud[37107]=16'hc077;
aud[37108]=16'hc074;
aud[37109]=16'hc072;
aud[37110]=16'hc06f;
aud[37111]=16'hc06d;
aud[37112]=16'hc06a;
aud[37113]=16'hc068;
aud[37114]=16'hc065;
aud[37115]=16'hc063;
aud[37116]=16'hc061;
aud[37117]=16'hc05e;
aud[37118]=16'hc05c;
aud[37119]=16'hc05a;
aud[37120]=16'hc058;
aud[37121]=16'hc055;
aud[37122]=16'hc053;
aud[37123]=16'hc051;
aud[37124]=16'hc04f;
aud[37125]=16'hc04d;
aud[37126]=16'hc04b;
aud[37127]=16'hc049;
aud[37128]=16'hc047;
aud[37129]=16'hc045;
aud[37130]=16'hc043;
aud[37131]=16'hc041;
aud[37132]=16'hc03f;
aud[37133]=16'hc03d;
aud[37134]=16'hc03b;
aud[37135]=16'hc039;
aud[37136]=16'hc038;
aud[37137]=16'hc036;
aud[37138]=16'hc034;
aud[37139]=16'hc033;
aud[37140]=16'hc031;
aud[37141]=16'hc02f;
aud[37142]=16'hc02e;
aud[37143]=16'hc02c;
aud[37144]=16'hc02a;
aud[37145]=16'hc029;
aud[37146]=16'hc027;
aud[37147]=16'hc026;
aud[37148]=16'hc024;
aud[37149]=16'hc023;
aud[37150]=16'hc022;
aud[37151]=16'hc020;
aud[37152]=16'hc01f;
aud[37153]=16'hc01e;
aud[37154]=16'hc01c;
aud[37155]=16'hc01b;
aud[37156]=16'hc01a;
aud[37157]=16'hc019;
aud[37158]=16'hc018;
aud[37159]=16'hc016;
aud[37160]=16'hc015;
aud[37161]=16'hc014;
aud[37162]=16'hc013;
aud[37163]=16'hc012;
aud[37164]=16'hc011;
aud[37165]=16'hc010;
aud[37166]=16'hc00f;
aud[37167]=16'hc00e;
aud[37168]=16'hc00d;
aud[37169]=16'hc00d;
aud[37170]=16'hc00c;
aud[37171]=16'hc00b;
aud[37172]=16'hc00a;
aud[37173]=16'hc009;
aud[37174]=16'hc009;
aud[37175]=16'hc008;
aud[37176]=16'hc007;
aud[37177]=16'hc007;
aud[37178]=16'hc006;
aud[37179]=16'hc006;
aud[37180]=16'hc005;
aud[37181]=16'hc005;
aud[37182]=16'hc004;
aud[37183]=16'hc004;
aud[37184]=16'hc003;
aud[37185]=16'hc003;
aud[37186]=16'hc002;
aud[37187]=16'hc002;
aud[37188]=16'hc002;
aud[37189]=16'hc001;
aud[37190]=16'hc001;
aud[37191]=16'hc001;
aud[37192]=16'hc001;
aud[37193]=16'hc001;
aud[37194]=16'hc000;
aud[37195]=16'hc000;
aud[37196]=16'hc000;
aud[37197]=16'hc000;
aud[37198]=16'hc000;
aud[37199]=16'hc000;
aud[37200]=16'hc000;
aud[37201]=16'hc000;
aud[37202]=16'hc000;
aud[37203]=16'hc000;
aud[37204]=16'hc000;
aud[37205]=16'hc001;
aud[37206]=16'hc001;
aud[37207]=16'hc001;
aud[37208]=16'hc001;
aud[37209]=16'hc001;
aud[37210]=16'hc002;
aud[37211]=16'hc002;
aud[37212]=16'hc002;
aud[37213]=16'hc003;
aud[37214]=16'hc003;
aud[37215]=16'hc004;
aud[37216]=16'hc004;
aud[37217]=16'hc005;
aud[37218]=16'hc005;
aud[37219]=16'hc006;
aud[37220]=16'hc006;
aud[37221]=16'hc007;
aud[37222]=16'hc007;
aud[37223]=16'hc008;
aud[37224]=16'hc009;
aud[37225]=16'hc009;
aud[37226]=16'hc00a;
aud[37227]=16'hc00b;
aud[37228]=16'hc00c;
aud[37229]=16'hc00d;
aud[37230]=16'hc00d;
aud[37231]=16'hc00e;
aud[37232]=16'hc00f;
aud[37233]=16'hc010;
aud[37234]=16'hc011;
aud[37235]=16'hc012;
aud[37236]=16'hc013;
aud[37237]=16'hc014;
aud[37238]=16'hc015;
aud[37239]=16'hc016;
aud[37240]=16'hc018;
aud[37241]=16'hc019;
aud[37242]=16'hc01a;
aud[37243]=16'hc01b;
aud[37244]=16'hc01c;
aud[37245]=16'hc01e;
aud[37246]=16'hc01f;
aud[37247]=16'hc020;
aud[37248]=16'hc022;
aud[37249]=16'hc023;
aud[37250]=16'hc024;
aud[37251]=16'hc026;
aud[37252]=16'hc027;
aud[37253]=16'hc029;
aud[37254]=16'hc02a;
aud[37255]=16'hc02c;
aud[37256]=16'hc02e;
aud[37257]=16'hc02f;
aud[37258]=16'hc031;
aud[37259]=16'hc033;
aud[37260]=16'hc034;
aud[37261]=16'hc036;
aud[37262]=16'hc038;
aud[37263]=16'hc039;
aud[37264]=16'hc03b;
aud[37265]=16'hc03d;
aud[37266]=16'hc03f;
aud[37267]=16'hc041;
aud[37268]=16'hc043;
aud[37269]=16'hc045;
aud[37270]=16'hc047;
aud[37271]=16'hc049;
aud[37272]=16'hc04b;
aud[37273]=16'hc04d;
aud[37274]=16'hc04f;
aud[37275]=16'hc051;
aud[37276]=16'hc053;
aud[37277]=16'hc055;
aud[37278]=16'hc058;
aud[37279]=16'hc05a;
aud[37280]=16'hc05c;
aud[37281]=16'hc05e;
aud[37282]=16'hc061;
aud[37283]=16'hc063;
aud[37284]=16'hc065;
aud[37285]=16'hc068;
aud[37286]=16'hc06a;
aud[37287]=16'hc06d;
aud[37288]=16'hc06f;
aud[37289]=16'hc072;
aud[37290]=16'hc074;
aud[37291]=16'hc077;
aud[37292]=16'hc079;
aud[37293]=16'hc07c;
aud[37294]=16'hc07f;
aud[37295]=16'hc081;
aud[37296]=16'hc084;
aud[37297]=16'hc087;
aud[37298]=16'hc089;
aud[37299]=16'hc08c;
aud[37300]=16'hc08f;
aud[37301]=16'hc092;
aud[37302]=16'hc095;
aud[37303]=16'hc098;
aud[37304]=16'hc09b;
aud[37305]=16'hc09d;
aud[37306]=16'hc0a0;
aud[37307]=16'hc0a3;
aud[37308]=16'hc0a6;
aud[37309]=16'hc0aa;
aud[37310]=16'hc0ad;
aud[37311]=16'hc0b0;
aud[37312]=16'hc0b3;
aud[37313]=16'hc0b6;
aud[37314]=16'hc0b9;
aud[37315]=16'hc0bd;
aud[37316]=16'hc0c0;
aud[37317]=16'hc0c3;
aud[37318]=16'hc0c6;
aud[37319]=16'hc0ca;
aud[37320]=16'hc0cd;
aud[37321]=16'hc0d0;
aud[37322]=16'hc0d4;
aud[37323]=16'hc0d7;
aud[37324]=16'hc0db;
aud[37325]=16'hc0de;
aud[37326]=16'hc0e2;
aud[37327]=16'hc0e5;
aud[37328]=16'hc0e9;
aud[37329]=16'hc0ed;
aud[37330]=16'hc0f0;
aud[37331]=16'hc0f4;
aud[37332]=16'hc0f8;
aud[37333]=16'hc0fb;
aud[37334]=16'hc0ff;
aud[37335]=16'hc103;
aud[37336]=16'hc107;
aud[37337]=16'hc10b;
aud[37338]=16'hc10e;
aud[37339]=16'hc112;
aud[37340]=16'hc116;
aud[37341]=16'hc11a;
aud[37342]=16'hc11e;
aud[37343]=16'hc122;
aud[37344]=16'hc126;
aud[37345]=16'hc12a;
aud[37346]=16'hc12e;
aud[37347]=16'hc133;
aud[37348]=16'hc137;
aud[37349]=16'hc13b;
aud[37350]=16'hc13f;
aud[37351]=16'hc143;
aud[37352]=16'hc147;
aud[37353]=16'hc14c;
aud[37354]=16'hc150;
aud[37355]=16'hc154;
aud[37356]=16'hc159;
aud[37357]=16'hc15d;
aud[37358]=16'hc162;
aud[37359]=16'hc166;
aud[37360]=16'hc16b;
aud[37361]=16'hc16f;
aud[37362]=16'hc174;
aud[37363]=16'hc178;
aud[37364]=16'hc17d;
aud[37365]=16'hc181;
aud[37366]=16'hc186;
aud[37367]=16'hc18b;
aud[37368]=16'hc18f;
aud[37369]=16'hc194;
aud[37370]=16'hc199;
aud[37371]=16'hc19e;
aud[37372]=16'hc1a2;
aud[37373]=16'hc1a7;
aud[37374]=16'hc1ac;
aud[37375]=16'hc1b1;
aud[37376]=16'hc1b6;
aud[37377]=16'hc1bb;
aud[37378]=16'hc1c0;
aud[37379]=16'hc1c5;
aud[37380]=16'hc1ca;
aud[37381]=16'hc1cf;
aud[37382]=16'hc1d4;
aud[37383]=16'hc1d9;
aud[37384]=16'hc1de;
aud[37385]=16'hc1e3;
aud[37386]=16'hc1e8;
aud[37387]=16'hc1ee;
aud[37388]=16'hc1f3;
aud[37389]=16'hc1f8;
aud[37390]=16'hc1fd;
aud[37391]=16'hc203;
aud[37392]=16'hc208;
aud[37393]=16'hc20d;
aud[37394]=16'hc213;
aud[37395]=16'hc218;
aud[37396]=16'hc21e;
aud[37397]=16'hc223;
aud[37398]=16'hc229;
aud[37399]=16'hc22e;
aud[37400]=16'hc234;
aud[37401]=16'hc239;
aud[37402]=16'hc23f;
aud[37403]=16'hc245;
aud[37404]=16'hc24a;
aud[37405]=16'hc250;
aud[37406]=16'hc256;
aud[37407]=16'hc25c;
aud[37408]=16'hc261;
aud[37409]=16'hc267;
aud[37410]=16'hc26d;
aud[37411]=16'hc273;
aud[37412]=16'hc279;
aud[37413]=16'hc27f;
aud[37414]=16'hc285;
aud[37415]=16'hc28b;
aud[37416]=16'hc291;
aud[37417]=16'hc297;
aud[37418]=16'hc29d;
aud[37419]=16'hc2a3;
aud[37420]=16'hc2a9;
aud[37421]=16'hc2af;
aud[37422]=16'hc2b5;
aud[37423]=16'hc2bb;
aud[37424]=16'hc2c1;
aud[37425]=16'hc2c8;
aud[37426]=16'hc2ce;
aud[37427]=16'hc2d4;
aud[37428]=16'hc2db;
aud[37429]=16'hc2e1;
aud[37430]=16'hc2e7;
aud[37431]=16'hc2ee;
aud[37432]=16'hc2f4;
aud[37433]=16'hc2fb;
aud[37434]=16'hc301;
aud[37435]=16'hc308;
aud[37436]=16'hc30e;
aud[37437]=16'hc315;
aud[37438]=16'hc31b;
aud[37439]=16'hc322;
aud[37440]=16'hc329;
aud[37441]=16'hc32f;
aud[37442]=16'hc336;
aud[37443]=16'hc33d;
aud[37444]=16'hc343;
aud[37445]=16'hc34a;
aud[37446]=16'hc351;
aud[37447]=16'hc358;
aud[37448]=16'hc35f;
aud[37449]=16'hc365;
aud[37450]=16'hc36c;
aud[37451]=16'hc373;
aud[37452]=16'hc37a;
aud[37453]=16'hc381;
aud[37454]=16'hc388;
aud[37455]=16'hc38f;
aud[37456]=16'hc396;
aud[37457]=16'hc39d;
aud[37458]=16'hc3a5;
aud[37459]=16'hc3ac;
aud[37460]=16'hc3b3;
aud[37461]=16'hc3ba;
aud[37462]=16'hc3c1;
aud[37463]=16'hc3c9;
aud[37464]=16'hc3d0;
aud[37465]=16'hc3d7;
aud[37466]=16'hc3df;
aud[37467]=16'hc3e6;
aud[37468]=16'hc3ed;
aud[37469]=16'hc3f5;
aud[37470]=16'hc3fc;
aud[37471]=16'hc404;
aud[37472]=16'hc40b;
aud[37473]=16'hc413;
aud[37474]=16'hc41a;
aud[37475]=16'hc422;
aud[37476]=16'hc429;
aud[37477]=16'hc431;
aud[37478]=16'hc439;
aud[37479]=16'hc440;
aud[37480]=16'hc448;
aud[37481]=16'hc450;
aud[37482]=16'hc457;
aud[37483]=16'hc45f;
aud[37484]=16'hc467;
aud[37485]=16'hc46f;
aud[37486]=16'hc477;
aud[37487]=16'hc47f;
aud[37488]=16'hc486;
aud[37489]=16'hc48e;
aud[37490]=16'hc496;
aud[37491]=16'hc49e;
aud[37492]=16'hc4a6;
aud[37493]=16'hc4ae;
aud[37494]=16'hc4b6;
aud[37495]=16'hc4bf;
aud[37496]=16'hc4c7;
aud[37497]=16'hc4cf;
aud[37498]=16'hc4d7;
aud[37499]=16'hc4df;
aud[37500]=16'hc4e7;
aud[37501]=16'hc4f0;
aud[37502]=16'hc4f8;
aud[37503]=16'hc500;
aud[37504]=16'hc509;
aud[37505]=16'hc511;
aud[37506]=16'hc519;
aud[37507]=16'hc522;
aud[37508]=16'hc52a;
aud[37509]=16'hc533;
aud[37510]=16'hc53b;
aud[37511]=16'hc544;
aud[37512]=16'hc54c;
aud[37513]=16'hc555;
aud[37514]=16'hc55d;
aud[37515]=16'hc566;
aud[37516]=16'hc56e;
aud[37517]=16'hc577;
aud[37518]=16'hc580;
aud[37519]=16'hc588;
aud[37520]=16'hc591;
aud[37521]=16'hc59a;
aud[37522]=16'hc5a3;
aud[37523]=16'hc5ac;
aud[37524]=16'hc5b4;
aud[37525]=16'hc5bd;
aud[37526]=16'hc5c6;
aud[37527]=16'hc5cf;
aud[37528]=16'hc5d8;
aud[37529]=16'hc5e1;
aud[37530]=16'hc5ea;
aud[37531]=16'hc5f3;
aud[37532]=16'hc5fc;
aud[37533]=16'hc605;
aud[37534]=16'hc60e;
aud[37535]=16'hc617;
aud[37536]=16'hc620;
aud[37537]=16'hc62a;
aud[37538]=16'hc633;
aud[37539]=16'hc63c;
aud[37540]=16'hc645;
aud[37541]=16'hc64f;
aud[37542]=16'hc658;
aud[37543]=16'hc661;
aud[37544]=16'hc66b;
aud[37545]=16'hc674;
aud[37546]=16'hc67d;
aud[37547]=16'hc687;
aud[37548]=16'hc690;
aud[37549]=16'hc69a;
aud[37550]=16'hc6a3;
aud[37551]=16'hc6ad;
aud[37552]=16'hc6b6;
aud[37553]=16'hc6c0;
aud[37554]=16'hc6c9;
aud[37555]=16'hc6d3;
aud[37556]=16'hc6dd;
aud[37557]=16'hc6e6;
aud[37558]=16'hc6f0;
aud[37559]=16'hc6fa;
aud[37560]=16'hc703;
aud[37561]=16'hc70d;
aud[37562]=16'hc717;
aud[37563]=16'hc721;
aud[37564]=16'hc72b;
aud[37565]=16'hc735;
aud[37566]=16'hc73f;
aud[37567]=16'hc748;
aud[37568]=16'hc752;
aud[37569]=16'hc75c;
aud[37570]=16'hc766;
aud[37571]=16'hc770;
aud[37572]=16'hc77a;
aud[37573]=16'hc785;
aud[37574]=16'hc78f;
aud[37575]=16'hc799;
aud[37576]=16'hc7a3;
aud[37577]=16'hc7ad;
aud[37578]=16'hc7b7;
aud[37579]=16'hc7c1;
aud[37580]=16'hc7cc;
aud[37581]=16'hc7d6;
aud[37582]=16'hc7e0;
aud[37583]=16'hc7eb;
aud[37584]=16'hc7f5;
aud[37585]=16'hc7ff;
aud[37586]=16'hc80a;
aud[37587]=16'hc814;
aud[37588]=16'hc81f;
aud[37589]=16'hc829;
aud[37590]=16'hc834;
aud[37591]=16'hc83e;
aud[37592]=16'hc849;
aud[37593]=16'hc853;
aud[37594]=16'hc85e;
aud[37595]=16'hc868;
aud[37596]=16'hc873;
aud[37597]=16'hc87e;
aud[37598]=16'hc888;
aud[37599]=16'hc893;
aud[37600]=16'hc89e;
aud[37601]=16'hc8a9;
aud[37602]=16'hc8b3;
aud[37603]=16'hc8be;
aud[37604]=16'hc8c9;
aud[37605]=16'hc8d4;
aud[37606]=16'hc8df;
aud[37607]=16'hc8ea;
aud[37608]=16'hc8f5;
aud[37609]=16'hc8ff;
aud[37610]=16'hc90a;
aud[37611]=16'hc915;
aud[37612]=16'hc920;
aud[37613]=16'hc92c;
aud[37614]=16'hc937;
aud[37615]=16'hc942;
aud[37616]=16'hc94d;
aud[37617]=16'hc958;
aud[37618]=16'hc963;
aud[37619]=16'hc96e;
aud[37620]=16'hc97a;
aud[37621]=16'hc985;
aud[37622]=16'hc990;
aud[37623]=16'hc99b;
aud[37624]=16'hc9a7;
aud[37625]=16'hc9b2;
aud[37626]=16'hc9bd;
aud[37627]=16'hc9c9;
aud[37628]=16'hc9d4;
aud[37629]=16'hc9e0;
aud[37630]=16'hc9eb;
aud[37631]=16'hc9f7;
aud[37632]=16'hca02;
aud[37633]=16'hca0e;
aud[37634]=16'hca19;
aud[37635]=16'hca25;
aud[37636]=16'hca30;
aud[37637]=16'hca3c;
aud[37638]=16'hca48;
aud[37639]=16'hca53;
aud[37640]=16'hca5f;
aud[37641]=16'hca6b;
aud[37642]=16'hca76;
aud[37643]=16'hca82;
aud[37644]=16'hca8e;
aud[37645]=16'hca9a;
aud[37646]=16'hcaa6;
aud[37647]=16'hcab1;
aud[37648]=16'hcabd;
aud[37649]=16'hcac9;
aud[37650]=16'hcad5;
aud[37651]=16'hcae1;
aud[37652]=16'hcaed;
aud[37653]=16'hcaf9;
aud[37654]=16'hcb05;
aud[37655]=16'hcb11;
aud[37656]=16'hcb1d;
aud[37657]=16'hcb29;
aud[37658]=16'hcb35;
aud[37659]=16'hcb42;
aud[37660]=16'hcb4e;
aud[37661]=16'hcb5a;
aud[37662]=16'hcb66;
aud[37663]=16'hcb72;
aud[37664]=16'hcb7f;
aud[37665]=16'hcb8b;
aud[37666]=16'hcb97;
aud[37667]=16'hcba3;
aud[37668]=16'hcbb0;
aud[37669]=16'hcbbc;
aud[37670]=16'hcbc9;
aud[37671]=16'hcbd5;
aud[37672]=16'hcbe1;
aud[37673]=16'hcbee;
aud[37674]=16'hcbfa;
aud[37675]=16'hcc07;
aud[37676]=16'hcc13;
aud[37677]=16'hcc20;
aud[37678]=16'hcc2c;
aud[37679]=16'hcc39;
aud[37680]=16'hcc46;
aud[37681]=16'hcc52;
aud[37682]=16'hcc5f;
aud[37683]=16'hcc6c;
aud[37684]=16'hcc78;
aud[37685]=16'hcc85;
aud[37686]=16'hcc92;
aud[37687]=16'hcc9f;
aud[37688]=16'hccab;
aud[37689]=16'hccb8;
aud[37690]=16'hccc5;
aud[37691]=16'hccd2;
aud[37692]=16'hccdf;
aud[37693]=16'hccec;
aud[37694]=16'hccf9;
aud[37695]=16'hcd06;
aud[37696]=16'hcd13;
aud[37697]=16'hcd20;
aud[37698]=16'hcd2d;
aud[37699]=16'hcd3a;
aud[37700]=16'hcd47;
aud[37701]=16'hcd54;
aud[37702]=16'hcd61;
aud[37703]=16'hcd6e;
aud[37704]=16'hcd7b;
aud[37705]=16'hcd88;
aud[37706]=16'hcd96;
aud[37707]=16'hcda3;
aud[37708]=16'hcdb0;
aud[37709]=16'hcdbd;
aud[37710]=16'hcdcb;
aud[37711]=16'hcdd8;
aud[37712]=16'hcde5;
aud[37713]=16'hcdf3;
aud[37714]=16'hce00;
aud[37715]=16'hce0d;
aud[37716]=16'hce1b;
aud[37717]=16'hce28;
aud[37718]=16'hce36;
aud[37719]=16'hce43;
aud[37720]=16'hce51;
aud[37721]=16'hce5e;
aud[37722]=16'hce6c;
aud[37723]=16'hce79;
aud[37724]=16'hce87;
aud[37725]=16'hce95;
aud[37726]=16'hcea2;
aud[37727]=16'hceb0;
aud[37728]=16'hcebe;
aud[37729]=16'hcecb;
aud[37730]=16'hced9;
aud[37731]=16'hcee7;
aud[37732]=16'hcef5;
aud[37733]=16'hcf02;
aud[37734]=16'hcf10;
aud[37735]=16'hcf1e;
aud[37736]=16'hcf2c;
aud[37737]=16'hcf3a;
aud[37738]=16'hcf48;
aud[37739]=16'hcf56;
aud[37740]=16'hcf63;
aud[37741]=16'hcf71;
aud[37742]=16'hcf7f;
aud[37743]=16'hcf8d;
aud[37744]=16'hcf9b;
aud[37745]=16'hcfa9;
aud[37746]=16'hcfb8;
aud[37747]=16'hcfc6;
aud[37748]=16'hcfd4;
aud[37749]=16'hcfe2;
aud[37750]=16'hcff0;
aud[37751]=16'hcffe;
aud[37752]=16'hd00c;
aud[37753]=16'hd01b;
aud[37754]=16'hd029;
aud[37755]=16'hd037;
aud[37756]=16'hd045;
aud[37757]=16'hd054;
aud[37758]=16'hd062;
aud[37759]=16'hd070;
aud[37760]=16'hd07f;
aud[37761]=16'hd08d;
aud[37762]=16'hd09b;
aud[37763]=16'hd0aa;
aud[37764]=16'hd0b8;
aud[37765]=16'hd0c7;
aud[37766]=16'hd0d5;
aud[37767]=16'hd0e4;
aud[37768]=16'hd0f2;
aud[37769]=16'hd101;
aud[37770]=16'hd10f;
aud[37771]=16'hd11e;
aud[37772]=16'hd12d;
aud[37773]=16'hd13b;
aud[37774]=16'hd14a;
aud[37775]=16'hd159;
aud[37776]=16'hd167;
aud[37777]=16'hd176;
aud[37778]=16'hd185;
aud[37779]=16'hd193;
aud[37780]=16'hd1a2;
aud[37781]=16'hd1b1;
aud[37782]=16'hd1c0;
aud[37783]=16'hd1cf;
aud[37784]=16'hd1de;
aud[37785]=16'hd1ec;
aud[37786]=16'hd1fb;
aud[37787]=16'hd20a;
aud[37788]=16'hd219;
aud[37789]=16'hd228;
aud[37790]=16'hd237;
aud[37791]=16'hd246;
aud[37792]=16'hd255;
aud[37793]=16'hd264;
aud[37794]=16'hd273;
aud[37795]=16'hd282;
aud[37796]=16'hd291;
aud[37797]=16'hd2a0;
aud[37798]=16'hd2b0;
aud[37799]=16'hd2bf;
aud[37800]=16'hd2ce;
aud[37801]=16'hd2dd;
aud[37802]=16'hd2ec;
aud[37803]=16'hd2fc;
aud[37804]=16'hd30b;
aud[37805]=16'hd31a;
aud[37806]=16'hd329;
aud[37807]=16'hd339;
aud[37808]=16'hd348;
aud[37809]=16'hd357;
aud[37810]=16'hd367;
aud[37811]=16'hd376;
aud[37812]=16'hd386;
aud[37813]=16'hd395;
aud[37814]=16'hd3a4;
aud[37815]=16'hd3b4;
aud[37816]=16'hd3c3;
aud[37817]=16'hd3d3;
aud[37818]=16'hd3e2;
aud[37819]=16'hd3f2;
aud[37820]=16'hd402;
aud[37821]=16'hd411;
aud[37822]=16'hd421;
aud[37823]=16'hd430;
aud[37824]=16'hd440;
aud[37825]=16'hd450;
aud[37826]=16'hd45f;
aud[37827]=16'hd46f;
aud[37828]=16'hd47f;
aud[37829]=16'hd48f;
aud[37830]=16'hd49e;
aud[37831]=16'hd4ae;
aud[37832]=16'hd4be;
aud[37833]=16'hd4ce;
aud[37834]=16'hd4de;
aud[37835]=16'hd4ed;
aud[37836]=16'hd4fd;
aud[37837]=16'hd50d;
aud[37838]=16'hd51d;
aud[37839]=16'hd52d;
aud[37840]=16'hd53d;
aud[37841]=16'hd54d;
aud[37842]=16'hd55d;
aud[37843]=16'hd56d;
aud[37844]=16'hd57d;
aud[37845]=16'hd58d;
aud[37846]=16'hd59d;
aud[37847]=16'hd5ad;
aud[37848]=16'hd5bd;
aud[37849]=16'hd5cd;
aud[37850]=16'hd5dd;
aud[37851]=16'hd5ee;
aud[37852]=16'hd5fe;
aud[37853]=16'hd60e;
aud[37854]=16'hd61e;
aud[37855]=16'hd62e;
aud[37856]=16'hd63f;
aud[37857]=16'hd64f;
aud[37858]=16'hd65f;
aud[37859]=16'hd66f;
aud[37860]=16'hd680;
aud[37861]=16'hd690;
aud[37862]=16'hd6a0;
aud[37863]=16'hd6b1;
aud[37864]=16'hd6c1;
aud[37865]=16'hd6d2;
aud[37866]=16'hd6e2;
aud[37867]=16'hd6f2;
aud[37868]=16'hd703;
aud[37869]=16'hd713;
aud[37870]=16'hd724;
aud[37871]=16'hd734;
aud[37872]=16'hd745;
aud[37873]=16'hd756;
aud[37874]=16'hd766;
aud[37875]=16'hd777;
aud[37876]=16'hd787;
aud[37877]=16'hd798;
aud[37878]=16'hd7a9;
aud[37879]=16'hd7b9;
aud[37880]=16'hd7ca;
aud[37881]=16'hd7db;
aud[37882]=16'hd7eb;
aud[37883]=16'hd7fc;
aud[37884]=16'hd80d;
aud[37885]=16'hd81e;
aud[37886]=16'hd82e;
aud[37887]=16'hd83f;
aud[37888]=16'hd850;
aud[37889]=16'hd861;
aud[37890]=16'hd872;
aud[37891]=16'hd882;
aud[37892]=16'hd893;
aud[37893]=16'hd8a4;
aud[37894]=16'hd8b5;
aud[37895]=16'hd8c6;
aud[37896]=16'hd8d7;
aud[37897]=16'hd8e8;
aud[37898]=16'hd8f9;
aud[37899]=16'hd90a;
aud[37900]=16'hd91b;
aud[37901]=16'hd92c;
aud[37902]=16'hd93d;
aud[37903]=16'hd94e;
aud[37904]=16'hd95f;
aud[37905]=16'hd970;
aud[37906]=16'hd982;
aud[37907]=16'hd993;
aud[37908]=16'hd9a4;
aud[37909]=16'hd9b5;
aud[37910]=16'hd9c6;
aud[37911]=16'hd9d7;
aud[37912]=16'hd9e9;
aud[37913]=16'hd9fa;
aud[37914]=16'hda0b;
aud[37915]=16'hda1c;
aud[37916]=16'hda2e;
aud[37917]=16'hda3f;
aud[37918]=16'hda50;
aud[37919]=16'hda62;
aud[37920]=16'hda73;
aud[37921]=16'hda84;
aud[37922]=16'hda96;
aud[37923]=16'hdaa7;
aud[37924]=16'hdab9;
aud[37925]=16'hdaca;
aud[37926]=16'hdadc;
aud[37927]=16'hdaed;
aud[37928]=16'hdaff;
aud[37929]=16'hdb10;
aud[37930]=16'hdb22;
aud[37931]=16'hdb33;
aud[37932]=16'hdb45;
aud[37933]=16'hdb56;
aud[37934]=16'hdb68;
aud[37935]=16'hdb79;
aud[37936]=16'hdb8b;
aud[37937]=16'hdb9d;
aud[37938]=16'hdbae;
aud[37939]=16'hdbc0;
aud[37940]=16'hdbd2;
aud[37941]=16'hdbe3;
aud[37942]=16'hdbf5;
aud[37943]=16'hdc07;
aud[37944]=16'hdc19;
aud[37945]=16'hdc2a;
aud[37946]=16'hdc3c;
aud[37947]=16'hdc4e;
aud[37948]=16'hdc60;
aud[37949]=16'hdc72;
aud[37950]=16'hdc83;
aud[37951]=16'hdc95;
aud[37952]=16'hdca7;
aud[37953]=16'hdcb9;
aud[37954]=16'hdccb;
aud[37955]=16'hdcdd;
aud[37956]=16'hdcef;
aud[37957]=16'hdd01;
aud[37958]=16'hdd13;
aud[37959]=16'hdd25;
aud[37960]=16'hdd37;
aud[37961]=16'hdd49;
aud[37962]=16'hdd5b;
aud[37963]=16'hdd6d;
aud[37964]=16'hdd7f;
aud[37965]=16'hdd91;
aud[37966]=16'hdda3;
aud[37967]=16'hddb5;
aud[37968]=16'hddc7;
aud[37969]=16'hddd9;
aud[37970]=16'hddeb;
aud[37971]=16'hddfe;
aud[37972]=16'hde10;
aud[37973]=16'hde22;
aud[37974]=16'hde34;
aud[37975]=16'hde46;
aud[37976]=16'hde59;
aud[37977]=16'hde6b;
aud[37978]=16'hde7d;
aud[37979]=16'hde8f;
aud[37980]=16'hdea2;
aud[37981]=16'hdeb4;
aud[37982]=16'hdec6;
aud[37983]=16'hded9;
aud[37984]=16'hdeeb;
aud[37985]=16'hdefd;
aud[37986]=16'hdf10;
aud[37987]=16'hdf22;
aud[37988]=16'hdf35;
aud[37989]=16'hdf47;
aud[37990]=16'hdf59;
aud[37991]=16'hdf6c;
aud[37992]=16'hdf7e;
aud[37993]=16'hdf91;
aud[37994]=16'hdfa3;
aud[37995]=16'hdfb6;
aud[37996]=16'hdfc8;
aud[37997]=16'hdfdb;
aud[37998]=16'hdfed;
aud[37999]=16'he000;
aud[38000]=16'he013;
aud[38001]=16'he025;
aud[38002]=16'he038;
aud[38003]=16'he04a;
aud[38004]=16'he05d;
aud[38005]=16'he070;
aud[38006]=16'he082;
aud[38007]=16'he095;
aud[38008]=16'he0a8;
aud[38009]=16'he0ba;
aud[38010]=16'he0cd;
aud[38011]=16'he0e0;
aud[38012]=16'he0f3;
aud[38013]=16'he105;
aud[38014]=16'he118;
aud[38015]=16'he12b;
aud[38016]=16'he13e;
aud[38017]=16'he151;
aud[38018]=16'he163;
aud[38019]=16'he176;
aud[38020]=16'he189;
aud[38021]=16'he19c;
aud[38022]=16'he1af;
aud[38023]=16'he1c2;
aud[38024]=16'he1d5;
aud[38025]=16'he1e8;
aud[38026]=16'he1fa;
aud[38027]=16'he20d;
aud[38028]=16'he220;
aud[38029]=16'he233;
aud[38030]=16'he246;
aud[38031]=16'he259;
aud[38032]=16'he26c;
aud[38033]=16'he27f;
aud[38034]=16'he292;
aud[38035]=16'he2a5;
aud[38036]=16'he2b9;
aud[38037]=16'he2cc;
aud[38038]=16'he2df;
aud[38039]=16'he2f2;
aud[38040]=16'he305;
aud[38041]=16'he318;
aud[38042]=16'he32b;
aud[38043]=16'he33e;
aud[38044]=16'he352;
aud[38045]=16'he365;
aud[38046]=16'he378;
aud[38047]=16'he38b;
aud[38048]=16'he39e;
aud[38049]=16'he3b2;
aud[38050]=16'he3c5;
aud[38051]=16'he3d8;
aud[38052]=16'he3eb;
aud[38053]=16'he3ff;
aud[38054]=16'he412;
aud[38055]=16'he425;
aud[38056]=16'he438;
aud[38057]=16'he44c;
aud[38058]=16'he45f;
aud[38059]=16'he473;
aud[38060]=16'he486;
aud[38061]=16'he499;
aud[38062]=16'he4ad;
aud[38063]=16'he4c0;
aud[38064]=16'he4d3;
aud[38065]=16'he4e7;
aud[38066]=16'he4fa;
aud[38067]=16'he50e;
aud[38068]=16'he521;
aud[38069]=16'he535;
aud[38070]=16'he548;
aud[38071]=16'he55c;
aud[38072]=16'he56f;
aud[38073]=16'he583;
aud[38074]=16'he596;
aud[38075]=16'he5aa;
aud[38076]=16'he5bd;
aud[38077]=16'he5d1;
aud[38078]=16'he5e4;
aud[38079]=16'he5f8;
aud[38080]=16'he60c;
aud[38081]=16'he61f;
aud[38082]=16'he633;
aud[38083]=16'he646;
aud[38084]=16'he65a;
aud[38085]=16'he66e;
aud[38086]=16'he681;
aud[38087]=16'he695;
aud[38088]=16'he6a9;
aud[38089]=16'he6bd;
aud[38090]=16'he6d0;
aud[38091]=16'he6e4;
aud[38092]=16'he6f8;
aud[38093]=16'he70b;
aud[38094]=16'he71f;
aud[38095]=16'he733;
aud[38096]=16'he747;
aud[38097]=16'he75b;
aud[38098]=16'he76e;
aud[38099]=16'he782;
aud[38100]=16'he796;
aud[38101]=16'he7aa;
aud[38102]=16'he7be;
aud[38103]=16'he7d1;
aud[38104]=16'he7e5;
aud[38105]=16'he7f9;
aud[38106]=16'he80d;
aud[38107]=16'he821;
aud[38108]=16'he835;
aud[38109]=16'he849;
aud[38110]=16'he85d;
aud[38111]=16'he871;
aud[38112]=16'he885;
aud[38113]=16'he899;
aud[38114]=16'he8ad;
aud[38115]=16'he8c0;
aud[38116]=16'he8d4;
aud[38117]=16'he8e8;
aud[38118]=16'he8fc;
aud[38119]=16'he910;
aud[38120]=16'he925;
aud[38121]=16'he939;
aud[38122]=16'he94d;
aud[38123]=16'he961;
aud[38124]=16'he975;
aud[38125]=16'he989;
aud[38126]=16'he99d;
aud[38127]=16'he9b1;
aud[38128]=16'he9c5;
aud[38129]=16'he9d9;
aud[38130]=16'he9ed;
aud[38131]=16'hea01;
aud[38132]=16'hea16;
aud[38133]=16'hea2a;
aud[38134]=16'hea3e;
aud[38135]=16'hea52;
aud[38136]=16'hea66;
aud[38137]=16'hea7a;
aud[38138]=16'hea8f;
aud[38139]=16'heaa3;
aud[38140]=16'heab7;
aud[38141]=16'heacb;
aud[38142]=16'heae0;
aud[38143]=16'heaf4;
aud[38144]=16'heb08;
aud[38145]=16'heb1c;
aud[38146]=16'heb31;
aud[38147]=16'heb45;
aud[38148]=16'heb59;
aud[38149]=16'heb6e;
aud[38150]=16'heb82;
aud[38151]=16'heb96;
aud[38152]=16'hebab;
aud[38153]=16'hebbf;
aud[38154]=16'hebd3;
aud[38155]=16'hebe8;
aud[38156]=16'hebfc;
aud[38157]=16'hec10;
aud[38158]=16'hec25;
aud[38159]=16'hec39;
aud[38160]=16'hec4d;
aud[38161]=16'hec62;
aud[38162]=16'hec76;
aud[38163]=16'hec8b;
aud[38164]=16'hec9f;
aud[38165]=16'hecb4;
aud[38166]=16'hecc8;
aud[38167]=16'hecdd;
aud[38168]=16'hecf1;
aud[38169]=16'hed05;
aud[38170]=16'hed1a;
aud[38171]=16'hed2e;
aud[38172]=16'hed43;
aud[38173]=16'hed57;
aud[38174]=16'hed6c;
aud[38175]=16'hed81;
aud[38176]=16'hed95;
aud[38177]=16'hedaa;
aud[38178]=16'hedbe;
aud[38179]=16'hedd3;
aud[38180]=16'hede7;
aud[38181]=16'hedfc;
aud[38182]=16'hee10;
aud[38183]=16'hee25;
aud[38184]=16'hee3a;
aud[38185]=16'hee4e;
aud[38186]=16'hee63;
aud[38187]=16'hee77;
aud[38188]=16'hee8c;
aud[38189]=16'heea1;
aud[38190]=16'heeb5;
aud[38191]=16'heeca;
aud[38192]=16'heedf;
aud[38193]=16'heef3;
aud[38194]=16'hef08;
aud[38195]=16'hef1d;
aud[38196]=16'hef31;
aud[38197]=16'hef46;
aud[38198]=16'hef5b;
aud[38199]=16'hef70;
aud[38200]=16'hef84;
aud[38201]=16'hef99;
aud[38202]=16'hefae;
aud[38203]=16'hefc2;
aud[38204]=16'hefd7;
aud[38205]=16'hefec;
aud[38206]=16'hf001;
aud[38207]=16'hf015;
aud[38208]=16'hf02a;
aud[38209]=16'hf03f;
aud[38210]=16'hf054;
aud[38211]=16'hf069;
aud[38212]=16'hf07d;
aud[38213]=16'hf092;
aud[38214]=16'hf0a7;
aud[38215]=16'hf0bc;
aud[38216]=16'hf0d1;
aud[38217]=16'hf0e6;
aud[38218]=16'hf0fa;
aud[38219]=16'hf10f;
aud[38220]=16'hf124;
aud[38221]=16'hf139;
aud[38222]=16'hf14e;
aud[38223]=16'hf163;
aud[38224]=16'hf178;
aud[38225]=16'hf18c;
aud[38226]=16'hf1a1;
aud[38227]=16'hf1b6;
aud[38228]=16'hf1cb;
aud[38229]=16'hf1e0;
aud[38230]=16'hf1f5;
aud[38231]=16'hf20a;
aud[38232]=16'hf21f;
aud[38233]=16'hf234;
aud[38234]=16'hf249;
aud[38235]=16'hf25e;
aud[38236]=16'hf273;
aud[38237]=16'hf288;
aud[38238]=16'hf29d;
aud[38239]=16'hf2b2;
aud[38240]=16'hf2c7;
aud[38241]=16'hf2dc;
aud[38242]=16'hf2f1;
aud[38243]=16'hf306;
aud[38244]=16'hf31b;
aud[38245]=16'hf330;
aud[38246]=16'hf345;
aud[38247]=16'hf35a;
aud[38248]=16'hf36f;
aud[38249]=16'hf384;
aud[38250]=16'hf399;
aud[38251]=16'hf3ae;
aud[38252]=16'hf3c3;
aud[38253]=16'hf3d8;
aud[38254]=16'hf3ed;
aud[38255]=16'hf402;
aud[38256]=16'hf417;
aud[38257]=16'hf42c;
aud[38258]=16'hf441;
aud[38259]=16'hf456;
aud[38260]=16'hf46b;
aud[38261]=16'hf480;
aud[38262]=16'hf496;
aud[38263]=16'hf4ab;
aud[38264]=16'hf4c0;
aud[38265]=16'hf4d5;
aud[38266]=16'hf4ea;
aud[38267]=16'hf4ff;
aud[38268]=16'hf514;
aud[38269]=16'hf529;
aud[38270]=16'hf53f;
aud[38271]=16'hf554;
aud[38272]=16'hf569;
aud[38273]=16'hf57e;
aud[38274]=16'hf593;
aud[38275]=16'hf5a8;
aud[38276]=16'hf5bd;
aud[38277]=16'hf5d3;
aud[38278]=16'hf5e8;
aud[38279]=16'hf5fd;
aud[38280]=16'hf612;
aud[38281]=16'hf627;
aud[38282]=16'hf63d;
aud[38283]=16'hf652;
aud[38284]=16'hf667;
aud[38285]=16'hf67c;
aud[38286]=16'hf691;
aud[38287]=16'hf6a7;
aud[38288]=16'hf6bc;
aud[38289]=16'hf6d1;
aud[38290]=16'hf6e6;
aud[38291]=16'hf6fb;
aud[38292]=16'hf711;
aud[38293]=16'hf726;
aud[38294]=16'hf73b;
aud[38295]=16'hf750;
aud[38296]=16'hf766;
aud[38297]=16'hf77b;
aud[38298]=16'hf790;
aud[38299]=16'hf7a5;
aud[38300]=16'hf7bb;
aud[38301]=16'hf7d0;
aud[38302]=16'hf7e5;
aud[38303]=16'hf7fb;
aud[38304]=16'hf810;
aud[38305]=16'hf825;
aud[38306]=16'hf83a;
aud[38307]=16'hf850;
aud[38308]=16'hf865;
aud[38309]=16'hf87a;
aud[38310]=16'hf890;
aud[38311]=16'hf8a5;
aud[38312]=16'hf8ba;
aud[38313]=16'hf8cf;
aud[38314]=16'hf8e5;
aud[38315]=16'hf8fa;
aud[38316]=16'hf90f;
aud[38317]=16'hf925;
aud[38318]=16'hf93a;
aud[38319]=16'hf94f;
aud[38320]=16'hf965;
aud[38321]=16'hf97a;
aud[38322]=16'hf98f;
aud[38323]=16'hf9a5;
aud[38324]=16'hf9ba;
aud[38325]=16'hf9cf;
aud[38326]=16'hf9e5;
aud[38327]=16'hf9fa;
aud[38328]=16'hfa0f;
aud[38329]=16'hfa25;
aud[38330]=16'hfa3a;
aud[38331]=16'hfa50;
aud[38332]=16'hfa65;
aud[38333]=16'hfa7a;
aud[38334]=16'hfa90;
aud[38335]=16'hfaa5;
aud[38336]=16'hfaba;
aud[38337]=16'hfad0;
aud[38338]=16'hfae5;
aud[38339]=16'hfafb;
aud[38340]=16'hfb10;
aud[38341]=16'hfb25;
aud[38342]=16'hfb3b;
aud[38343]=16'hfb50;
aud[38344]=16'hfb65;
aud[38345]=16'hfb7b;
aud[38346]=16'hfb90;
aud[38347]=16'hfba6;
aud[38348]=16'hfbbb;
aud[38349]=16'hfbd0;
aud[38350]=16'hfbe6;
aud[38351]=16'hfbfb;
aud[38352]=16'hfc11;
aud[38353]=16'hfc26;
aud[38354]=16'hfc3b;
aud[38355]=16'hfc51;
aud[38356]=16'hfc66;
aud[38357]=16'hfc7c;
aud[38358]=16'hfc91;
aud[38359]=16'hfca7;
aud[38360]=16'hfcbc;
aud[38361]=16'hfcd1;
aud[38362]=16'hfce7;
aud[38363]=16'hfcfc;
aud[38364]=16'hfd12;
aud[38365]=16'hfd27;
aud[38366]=16'hfd3c;
aud[38367]=16'hfd52;
aud[38368]=16'hfd67;
aud[38369]=16'hfd7d;
aud[38370]=16'hfd92;
aud[38371]=16'hfda8;
aud[38372]=16'hfdbd;
aud[38373]=16'hfdd2;
aud[38374]=16'hfde8;
aud[38375]=16'hfdfd;
aud[38376]=16'hfe13;
aud[38377]=16'hfe28;
aud[38378]=16'hfe3e;
aud[38379]=16'hfe53;
aud[38380]=16'hfe69;
aud[38381]=16'hfe7e;
aud[38382]=16'hfe93;
aud[38383]=16'hfea9;
aud[38384]=16'hfebe;
aud[38385]=16'hfed4;
aud[38386]=16'hfee9;
aud[38387]=16'hfeff;
aud[38388]=16'hff14;
aud[38389]=16'hff2a;
aud[38390]=16'hff3f;
aud[38391]=16'hff54;
aud[38392]=16'hff6a;
aud[38393]=16'hff7f;
aud[38394]=16'hff95;
aud[38395]=16'hffaa;
aud[38396]=16'hffc0;
aud[38397]=16'hffd5;
aud[38398]=16'hffeb;
aud[38399]=16'h0;
aud[38400]=16'h15;
aud[38401]=16'h2b;
aud[38402]=16'h40;
aud[38403]=16'h56;
aud[38404]=16'h6b;
aud[38405]=16'h81;
aud[38406]=16'h96;
aud[38407]=16'hac;
aud[38408]=16'hc1;
aud[38409]=16'hd6;
aud[38410]=16'hec;
aud[38411]=16'h101;
aud[38412]=16'h117;
aud[38413]=16'h12c;
aud[38414]=16'h142;
aud[38415]=16'h157;
aud[38416]=16'h16d;
aud[38417]=16'h182;
aud[38418]=16'h197;
aud[38419]=16'h1ad;
aud[38420]=16'h1c2;
aud[38421]=16'h1d8;
aud[38422]=16'h1ed;
aud[38423]=16'h203;
aud[38424]=16'h218;
aud[38425]=16'h22e;
aud[38426]=16'h243;
aud[38427]=16'h258;
aud[38428]=16'h26e;
aud[38429]=16'h283;
aud[38430]=16'h299;
aud[38431]=16'h2ae;
aud[38432]=16'h2c4;
aud[38433]=16'h2d9;
aud[38434]=16'h2ee;
aud[38435]=16'h304;
aud[38436]=16'h319;
aud[38437]=16'h32f;
aud[38438]=16'h344;
aud[38439]=16'h359;
aud[38440]=16'h36f;
aud[38441]=16'h384;
aud[38442]=16'h39a;
aud[38443]=16'h3af;
aud[38444]=16'h3c5;
aud[38445]=16'h3da;
aud[38446]=16'h3ef;
aud[38447]=16'h405;
aud[38448]=16'h41a;
aud[38449]=16'h430;
aud[38450]=16'h445;
aud[38451]=16'h45a;
aud[38452]=16'h470;
aud[38453]=16'h485;
aud[38454]=16'h49b;
aud[38455]=16'h4b0;
aud[38456]=16'h4c5;
aud[38457]=16'h4db;
aud[38458]=16'h4f0;
aud[38459]=16'h505;
aud[38460]=16'h51b;
aud[38461]=16'h530;
aud[38462]=16'h546;
aud[38463]=16'h55b;
aud[38464]=16'h570;
aud[38465]=16'h586;
aud[38466]=16'h59b;
aud[38467]=16'h5b0;
aud[38468]=16'h5c6;
aud[38469]=16'h5db;
aud[38470]=16'h5f1;
aud[38471]=16'h606;
aud[38472]=16'h61b;
aud[38473]=16'h631;
aud[38474]=16'h646;
aud[38475]=16'h65b;
aud[38476]=16'h671;
aud[38477]=16'h686;
aud[38478]=16'h69b;
aud[38479]=16'h6b1;
aud[38480]=16'h6c6;
aud[38481]=16'h6db;
aud[38482]=16'h6f1;
aud[38483]=16'h706;
aud[38484]=16'h71b;
aud[38485]=16'h731;
aud[38486]=16'h746;
aud[38487]=16'h75b;
aud[38488]=16'h770;
aud[38489]=16'h786;
aud[38490]=16'h79b;
aud[38491]=16'h7b0;
aud[38492]=16'h7c6;
aud[38493]=16'h7db;
aud[38494]=16'h7f0;
aud[38495]=16'h805;
aud[38496]=16'h81b;
aud[38497]=16'h830;
aud[38498]=16'h845;
aud[38499]=16'h85b;
aud[38500]=16'h870;
aud[38501]=16'h885;
aud[38502]=16'h89a;
aud[38503]=16'h8b0;
aud[38504]=16'h8c5;
aud[38505]=16'h8da;
aud[38506]=16'h8ef;
aud[38507]=16'h905;
aud[38508]=16'h91a;
aud[38509]=16'h92f;
aud[38510]=16'h944;
aud[38511]=16'h959;
aud[38512]=16'h96f;
aud[38513]=16'h984;
aud[38514]=16'h999;
aud[38515]=16'h9ae;
aud[38516]=16'h9c3;
aud[38517]=16'h9d9;
aud[38518]=16'h9ee;
aud[38519]=16'ha03;
aud[38520]=16'ha18;
aud[38521]=16'ha2d;
aud[38522]=16'ha43;
aud[38523]=16'ha58;
aud[38524]=16'ha6d;
aud[38525]=16'ha82;
aud[38526]=16'ha97;
aud[38527]=16'haac;
aud[38528]=16'hac1;
aud[38529]=16'had7;
aud[38530]=16'haec;
aud[38531]=16'hb01;
aud[38532]=16'hb16;
aud[38533]=16'hb2b;
aud[38534]=16'hb40;
aud[38535]=16'hb55;
aud[38536]=16'hb6a;
aud[38537]=16'hb80;
aud[38538]=16'hb95;
aud[38539]=16'hbaa;
aud[38540]=16'hbbf;
aud[38541]=16'hbd4;
aud[38542]=16'hbe9;
aud[38543]=16'hbfe;
aud[38544]=16'hc13;
aud[38545]=16'hc28;
aud[38546]=16'hc3d;
aud[38547]=16'hc52;
aud[38548]=16'hc67;
aud[38549]=16'hc7c;
aud[38550]=16'hc91;
aud[38551]=16'hca6;
aud[38552]=16'hcbb;
aud[38553]=16'hcd0;
aud[38554]=16'hce5;
aud[38555]=16'hcfa;
aud[38556]=16'hd0f;
aud[38557]=16'hd24;
aud[38558]=16'hd39;
aud[38559]=16'hd4e;
aud[38560]=16'hd63;
aud[38561]=16'hd78;
aud[38562]=16'hd8d;
aud[38563]=16'hda2;
aud[38564]=16'hdb7;
aud[38565]=16'hdcc;
aud[38566]=16'hde1;
aud[38567]=16'hdf6;
aud[38568]=16'he0b;
aud[38569]=16'he20;
aud[38570]=16'he35;
aud[38571]=16'he4a;
aud[38572]=16'he5f;
aud[38573]=16'he74;
aud[38574]=16'he88;
aud[38575]=16'he9d;
aud[38576]=16'heb2;
aud[38577]=16'hec7;
aud[38578]=16'hedc;
aud[38579]=16'hef1;
aud[38580]=16'hf06;
aud[38581]=16'hf1a;
aud[38582]=16'hf2f;
aud[38583]=16'hf44;
aud[38584]=16'hf59;
aud[38585]=16'hf6e;
aud[38586]=16'hf83;
aud[38587]=16'hf97;
aud[38588]=16'hfac;
aud[38589]=16'hfc1;
aud[38590]=16'hfd6;
aud[38591]=16'hfeb;
aud[38592]=16'hfff;
aud[38593]=16'h1014;
aud[38594]=16'h1029;
aud[38595]=16'h103e;
aud[38596]=16'h1052;
aud[38597]=16'h1067;
aud[38598]=16'h107c;
aud[38599]=16'h1090;
aud[38600]=16'h10a5;
aud[38601]=16'h10ba;
aud[38602]=16'h10cf;
aud[38603]=16'h10e3;
aud[38604]=16'h10f8;
aud[38605]=16'h110d;
aud[38606]=16'h1121;
aud[38607]=16'h1136;
aud[38608]=16'h114b;
aud[38609]=16'h115f;
aud[38610]=16'h1174;
aud[38611]=16'h1189;
aud[38612]=16'h119d;
aud[38613]=16'h11b2;
aud[38614]=16'h11c6;
aud[38615]=16'h11db;
aud[38616]=16'h11f0;
aud[38617]=16'h1204;
aud[38618]=16'h1219;
aud[38619]=16'h122d;
aud[38620]=16'h1242;
aud[38621]=16'h1256;
aud[38622]=16'h126b;
aud[38623]=16'h127f;
aud[38624]=16'h1294;
aud[38625]=16'h12a9;
aud[38626]=16'h12bd;
aud[38627]=16'h12d2;
aud[38628]=16'h12e6;
aud[38629]=16'h12fb;
aud[38630]=16'h130f;
aud[38631]=16'h1323;
aud[38632]=16'h1338;
aud[38633]=16'h134c;
aud[38634]=16'h1361;
aud[38635]=16'h1375;
aud[38636]=16'h138a;
aud[38637]=16'h139e;
aud[38638]=16'h13b3;
aud[38639]=16'h13c7;
aud[38640]=16'h13db;
aud[38641]=16'h13f0;
aud[38642]=16'h1404;
aud[38643]=16'h1418;
aud[38644]=16'h142d;
aud[38645]=16'h1441;
aud[38646]=16'h1455;
aud[38647]=16'h146a;
aud[38648]=16'h147e;
aud[38649]=16'h1492;
aud[38650]=16'h14a7;
aud[38651]=16'h14bb;
aud[38652]=16'h14cf;
aud[38653]=16'h14e4;
aud[38654]=16'h14f8;
aud[38655]=16'h150c;
aud[38656]=16'h1520;
aud[38657]=16'h1535;
aud[38658]=16'h1549;
aud[38659]=16'h155d;
aud[38660]=16'h1571;
aud[38661]=16'h1586;
aud[38662]=16'h159a;
aud[38663]=16'h15ae;
aud[38664]=16'h15c2;
aud[38665]=16'h15d6;
aud[38666]=16'h15ea;
aud[38667]=16'h15ff;
aud[38668]=16'h1613;
aud[38669]=16'h1627;
aud[38670]=16'h163b;
aud[38671]=16'h164f;
aud[38672]=16'h1663;
aud[38673]=16'h1677;
aud[38674]=16'h168b;
aud[38675]=16'h169f;
aud[38676]=16'h16b3;
aud[38677]=16'h16c7;
aud[38678]=16'h16db;
aud[38679]=16'h16f0;
aud[38680]=16'h1704;
aud[38681]=16'h1718;
aud[38682]=16'h172c;
aud[38683]=16'h1740;
aud[38684]=16'h1753;
aud[38685]=16'h1767;
aud[38686]=16'h177b;
aud[38687]=16'h178f;
aud[38688]=16'h17a3;
aud[38689]=16'h17b7;
aud[38690]=16'h17cb;
aud[38691]=16'h17df;
aud[38692]=16'h17f3;
aud[38693]=16'h1807;
aud[38694]=16'h181b;
aud[38695]=16'h182f;
aud[38696]=16'h1842;
aud[38697]=16'h1856;
aud[38698]=16'h186a;
aud[38699]=16'h187e;
aud[38700]=16'h1892;
aud[38701]=16'h18a5;
aud[38702]=16'h18b9;
aud[38703]=16'h18cd;
aud[38704]=16'h18e1;
aud[38705]=16'h18f5;
aud[38706]=16'h1908;
aud[38707]=16'h191c;
aud[38708]=16'h1930;
aud[38709]=16'h1943;
aud[38710]=16'h1957;
aud[38711]=16'h196b;
aud[38712]=16'h197f;
aud[38713]=16'h1992;
aud[38714]=16'h19a6;
aud[38715]=16'h19ba;
aud[38716]=16'h19cd;
aud[38717]=16'h19e1;
aud[38718]=16'h19f4;
aud[38719]=16'h1a08;
aud[38720]=16'h1a1c;
aud[38721]=16'h1a2f;
aud[38722]=16'h1a43;
aud[38723]=16'h1a56;
aud[38724]=16'h1a6a;
aud[38725]=16'h1a7d;
aud[38726]=16'h1a91;
aud[38727]=16'h1aa4;
aud[38728]=16'h1ab8;
aud[38729]=16'h1acb;
aud[38730]=16'h1adf;
aud[38731]=16'h1af2;
aud[38732]=16'h1b06;
aud[38733]=16'h1b19;
aud[38734]=16'h1b2d;
aud[38735]=16'h1b40;
aud[38736]=16'h1b53;
aud[38737]=16'h1b67;
aud[38738]=16'h1b7a;
aud[38739]=16'h1b8d;
aud[38740]=16'h1ba1;
aud[38741]=16'h1bb4;
aud[38742]=16'h1bc8;
aud[38743]=16'h1bdb;
aud[38744]=16'h1bee;
aud[38745]=16'h1c01;
aud[38746]=16'h1c15;
aud[38747]=16'h1c28;
aud[38748]=16'h1c3b;
aud[38749]=16'h1c4e;
aud[38750]=16'h1c62;
aud[38751]=16'h1c75;
aud[38752]=16'h1c88;
aud[38753]=16'h1c9b;
aud[38754]=16'h1cae;
aud[38755]=16'h1cc2;
aud[38756]=16'h1cd5;
aud[38757]=16'h1ce8;
aud[38758]=16'h1cfb;
aud[38759]=16'h1d0e;
aud[38760]=16'h1d21;
aud[38761]=16'h1d34;
aud[38762]=16'h1d47;
aud[38763]=16'h1d5b;
aud[38764]=16'h1d6e;
aud[38765]=16'h1d81;
aud[38766]=16'h1d94;
aud[38767]=16'h1da7;
aud[38768]=16'h1dba;
aud[38769]=16'h1dcd;
aud[38770]=16'h1de0;
aud[38771]=16'h1df3;
aud[38772]=16'h1e06;
aud[38773]=16'h1e18;
aud[38774]=16'h1e2b;
aud[38775]=16'h1e3e;
aud[38776]=16'h1e51;
aud[38777]=16'h1e64;
aud[38778]=16'h1e77;
aud[38779]=16'h1e8a;
aud[38780]=16'h1e9d;
aud[38781]=16'h1eaf;
aud[38782]=16'h1ec2;
aud[38783]=16'h1ed5;
aud[38784]=16'h1ee8;
aud[38785]=16'h1efb;
aud[38786]=16'h1f0d;
aud[38787]=16'h1f20;
aud[38788]=16'h1f33;
aud[38789]=16'h1f46;
aud[38790]=16'h1f58;
aud[38791]=16'h1f6b;
aud[38792]=16'h1f7e;
aud[38793]=16'h1f90;
aud[38794]=16'h1fa3;
aud[38795]=16'h1fb6;
aud[38796]=16'h1fc8;
aud[38797]=16'h1fdb;
aud[38798]=16'h1fed;
aud[38799]=16'h2000;
aud[38800]=16'h2013;
aud[38801]=16'h2025;
aud[38802]=16'h2038;
aud[38803]=16'h204a;
aud[38804]=16'h205d;
aud[38805]=16'h206f;
aud[38806]=16'h2082;
aud[38807]=16'h2094;
aud[38808]=16'h20a7;
aud[38809]=16'h20b9;
aud[38810]=16'h20cb;
aud[38811]=16'h20de;
aud[38812]=16'h20f0;
aud[38813]=16'h2103;
aud[38814]=16'h2115;
aud[38815]=16'h2127;
aud[38816]=16'h213a;
aud[38817]=16'h214c;
aud[38818]=16'h215e;
aud[38819]=16'h2171;
aud[38820]=16'h2183;
aud[38821]=16'h2195;
aud[38822]=16'h21a7;
aud[38823]=16'h21ba;
aud[38824]=16'h21cc;
aud[38825]=16'h21de;
aud[38826]=16'h21f0;
aud[38827]=16'h2202;
aud[38828]=16'h2215;
aud[38829]=16'h2227;
aud[38830]=16'h2239;
aud[38831]=16'h224b;
aud[38832]=16'h225d;
aud[38833]=16'h226f;
aud[38834]=16'h2281;
aud[38835]=16'h2293;
aud[38836]=16'h22a5;
aud[38837]=16'h22b7;
aud[38838]=16'h22c9;
aud[38839]=16'h22db;
aud[38840]=16'h22ed;
aud[38841]=16'h22ff;
aud[38842]=16'h2311;
aud[38843]=16'h2323;
aud[38844]=16'h2335;
aud[38845]=16'h2347;
aud[38846]=16'h2359;
aud[38847]=16'h236b;
aud[38848]=16'h237d;
aud[38849]=16'h238e;
aud[38850]=16'h23a0;
aud[38851]=16'h23b2;
aud[38852]=16'h23c4;
aud[38853]=16'h23d6;
aud[38854]=16'h23e7;
aud[38855]=16'h23f9;
aud[38856]=16'h240b;
aud[38857]=16'h241d;
aud[38858]=16'h242e;
aud[38859]=16'h2440;
aud[38860]=16'h2452;
aud[38861]=16'h2463;
aud[38862]=16'h2475;
aud[38863]=16'h2487;
aud[38864]=16'h2498;
aud[38865]=16'h24aa;
aud[38866]=16'h24bb;
aud[38867]=16'h24cd;
aud[38868]=16'h24de;
aud[38869]=16'h24f0;
aud[38870]=16'h2501;
aud[38871]=16'h2513;
aud[38872]=16'h2524;
aud[38873]=16'h2536;
aud[38874]=16'h2547;
aud[38875]=16'h2559;
aud[38876]=16'h256a;
aud[38877]=16'h257c;
aud[38878]=16'h258d;
aud[38879]=16'h259e;
aud[38880]=16'h25b0;
aud[38881]=16'h25c1;
aud[38882]=16'h25d2;
aud[38883]=16'h25e4;
aud[38884]=16'h25f5;
aud[38885]=16'h2606;
aud[38886]=16'h2617;
aud[38887]=16'h2629;
aud[38888]=16'h263a;
aud[38889]=16'h264b;
aud[38890]=16'h265c;
aud[38891]=16'h266d;
aud[38892]=16'h267e;
aud[38893]=16'h2690;
aud[38894]=16'h26a1;
aud[38895]=16'h26b2;
aud[38896]=16'h26c3;
aud[38897]=16'h26d4;
aud[38898]=16'h26e5;
aud[38899]=16'h26f6;
aud[38900]=16'h2707;
aud[38901]=16'h2718;
aud[38902]=16'h2729;
aud[38903]=16'h273a;
aud[38904]=16'h274b;
aud[38905]=16'h275c;
aud[38906]=16'h276d;
aud[38907]=16'h277e;
aud[38908]=16'h278e;
aud[38909]=16'h279f;
aud[38910]=16'h27b0;
aud[38911]=16'h27c1;
aud[38912]=16'h27d2;
aud[38913]=16'h27e2;
aud[38914]=16'h27f3;
aud[38915]=16'h2804;
aud[38916]=16'h2815;
aud[38917]=16'h2825;
aud[38918]=16'h2836;
aud[38919]=16'h2847;
aud[38920]=16'h2857;
aud[38921]=16'h2868;
aud[38922]=16'h2879;
aud[38923]=16'h2889;
aud[38924]=16'h289a;
aud[38925]=16'h28aa;
aud[38926]=16'h28bb;
aud[38927]=16'h28cc;
aud[38928]=16'h28dc;
aud[38929]=16'h28ed;
aud[38930]=16'h28fd;
aud[38931]=16'h290e;
aud[38932]=16'h291e;
aud[38933]=16'h292e;
aud[38934]=16'h293f;
aud[38935]=16'h294f;
aud[38936]=16'h2960;
aud[38937]=16'h2970;
aud[38938]=16'h2980;
aud[38939]=16'h2991;
aud[38940]=16'h29a1;
aud[38941]=16'h29b1;
aud[38942]=16'h29c1;
aud[38943]=16'h29d2;
aud[38944]=16'h29e2;
aud[38945]=16'h29f2;
aud[38946]=16'h2a02;
aud[38947]=16'h2a12;
aud[38948]=16'h2a23;
aud[38949]=16'h2a33;
aud[38950]=16'h2a43;
aud[38951]=16'h2a53;
aud[38952]=16'h2a63;
aud[38953]=16'h2a73;
aud[38954]=16'h2a83;
aud[38955]=16'h2a93;
aud[38956]=16'h2aa3;
aud[38957]=16'h2ab3;
aud[38958]=16'h2ac3;
aud[38959]=16'h2ad3;
aud[38960]=16'h2ae3;
aud[38961]=16'h2af3;
aud[38962]=16'h2b03;
aud[38963]=16'h2b13;
aud[38964]=16'h2b22;
aud[38965]=16'h2b32;
aud[38966]=16'h2b42;
aud[38967]=16'h2b52;
aud[38968]=16'h2b62;
aud[38969]=16'h2b71;
aud[38970]=16'h2b81;
aud[38971]=16'h2b91;
aud[38972]=16'h2ba1;
aud[38973]=16'h2bb0;
aud[38974]=16'h2bc0;
aud[38975]=16'h2bd0;
aud[38976]=16'h2bdf;
aud[38977]=16'h2bef;
aud[38978]=16'h2bfe;
aud[38979]=16'h2c0e;
aud[38980]=16'h2c1e;
aud[38981]=16'h2c2d;
aud[38982]=16'h2c3d;
aud[38983]=16'h2c4c;
aud[38984]=16'h2c5c;
aud[38985]=16'h2c6b;
aud[38986]=16'h2c7a;
aud[38987]=16'h2c8a;
aud[38988]=16'h2c99;
aud[38989]=16'h2ca9;
aud[38990]=16'h2cb8;
aud[38991]=16'h2cc7;
aud[38992]=16'h2cd7;
aud[38993]=16'h2ce6;
aud[38994]=16'h2cf5;
aud[38995]=16'h2d04;
aud[38996]=16'h2d14;
aud[38997]=16'h2d23;
aud[38998]=16'h2d32;
aud[38999]=16'h2d41;
aud[39000]=16'h2d50;
aud[39001]=16'h2d60;
aud[39002]=16'h2d6f;
aud[39003]=16'h2d7e;
aud[39004]=16'h2d8d;
aud[39005]=16'h2d9c;
aud[39006]=16'h2dab;
aud[39007]=16'h2dba;
aud[39008]=16'h2dc9;
aud[39009]=16'h2dd8;
aud[39010]=16'h2de7;
aud[39011]=16'h2df6;
aud[39012]=16'h2e05;
aud[39013]=16'h2e14;
aud[39014]=16'h2e22;
aud[39015]=16'h2e31;
aud[39016]=16'h2e40;
aud[39017]=16'h2e4f;
aud[39018]=16'h2e5e;
aud[39019]=16'h2e6d;
aud[39020]=16'h2e7b;
aud[39021]=16'h2e8a;
aud[39022]=16'h2e99;
aud[39023]=16'h2ea7;
aud[39024]=16'h2eb6;
aud[39025]=16'h2ec5;
aud[39026]=16'h2ed3;
aud[39027]=16'h2ee2;
aud[39028]=16'h2ef1;
aud[39029]=16'h2eff;
aud[39030]=16'h2f0e;
aud[39031]=16'h2f1c;
aud[39032]=16'h2f2b;
aud[39033]=16'h2f39;
aud[39034]=16'h2f48;
aud[39035]=16'h2f56;
aud[39036]=16'h2f65;
aud[39037]=16'h2f73;
aud[39038]=16'h2f81;
aud[39039]=16'h2f90;
aud[39040]=16'h2f9e;
aud[39041]=16'h2fac;
aud[39042]=16'h2fbb;
aud[39043]=16'h2fc9;
aud[39044]=16'h2fd7;
aud[39045]=16'h2fe5;
aud[39046]=16'h2ff4;
aud[39047]=16'h3002;
aud[39048]=16'h3010;
aud[39049]=16'h301e;
aud[39050]=16'h302c;
aud[39051]=16'h303a;
aud[39052]=16'h3048;
aud[39053]=16'h3057;
aud[39054]=16'h3065;
aud[39055]=16'h3073;
aud[39056]=16'h3081;
aud[39057]=16'h308f;
aud[39058]=16'h309d;
aud[39059]=16'h30aa;
aud[39060]=16'h30b8;
aud[39061]=16'h30c6;
aud[39062]=16'h30d4;
aud[39063]=16'h30e2;
aud[39064]=16'h30f0;
aud[39065]=16'h30fe;
aud[39066]=16'h310b;
aud[39067]=16'h3119;
aud[39068]=16'h3127;
aud[39069]=16'h3135;
aud[39070]=16'h3142;
aud[39071]=16'h3150;
aud[39072]=16'h315e;
aud[39073]=16'h316b;
aud[39074]=16'h3179;
aud[39075]=16'h3187;
aud[39076]=16'h3194;
aud[39077]=16'h31a2;
aud[39078]=16'h31af;
aud[39079]=16'h31bd;
aud[39080]=16'h31ca;
aud[39081]=16'h31d8;
aud[39082]=16'h31e5;
aud[39083]=16'h31f3;
aud[39084]=16'h3200;
aud[39085]=16'h320d;
aud[39086]=16'h321b;
aud[39087]=16'h3228;
aud[39088]=16'h3235;
aud[39089]=16'h3243;
aud[39090]=16'h3250;
aud[39091]=16'h325d;
aud[39092]=16'h326a;
aud[39093]=16'h3278;
aud[39094]=16'h3285;
aud[39095]=16'h3292;
aud[39096]=16'h329f;
aud[39097]=16'h32ac;
aud[39098]=16'h32b9;
aud[39099]=16'h32c6;
aud[39100]=16'h32d3;
aud[39101]=16'h32e0;
aud[39102]=16'h32ed;
aud[39103]=16'h32fa;
aud[39104]=16'h3307;
aud[39105]=16'h3314;
aud[39106]=16'h3321;
aud[39107]=16'h332e;
aud[39108]=16'h333b;
aud[39109]=16'h3348;
aud[39110]=16'h3355;
aud[39111]=16'h3361;
aud[39112]=16'h336e;
aud[39113]=16'h337b;
aud[39114]=16'h3388;
aud[39115]=16'h3394;
aud[39116]=16'h33a1;
aud[39117]=16'h33ae;
aud[39118]=16'h33ba;
aud[39119]=16'h33c7;
aud[39120]=16'h33d4;
aud[39121]=16'h33e0;
aud[39122]=16'h33ed;
aud[39123]=16'h33f9;
aud[39124]=16'h3406;
aud[39125]=16'h3412;
aud[39126]=16'h341f;
aud[39127]=16'h342b;
aud[39128]=16'h3437;
aud[39129]=16'h3444;
aud[39130]=16'h3450;
aud[39131]=16'h345d;
aud[39132]=16'h3469;
aud[39133]=16'h3475;
aud[39134]=16'h3481;
aud[39135]=16'h348e;
aud[39136]=16'h349a;
aud[39137]=16'h34a6;
aud[39138]=16'h34b2;
aud[39139]=16'h34be;
aud[39140]=16'h34cb;
aud[39141]=16'h34d7;
aud[39142]=16'h34e3;
aud[39143]=16'h34ef;
aud[39144]=16'h34fb;
aud[39145]=16'h3507;
aud[39146]=16'h3513;
aud[39147]=16'h351f;
aud[39148]=16'h352b;
aud[39149]=16'h3537;
aud[39150]=16'h3543;
aud[39151]=16'h354f;
aud[39152]=16'h355a;
aud[39153]=16'h3566;
aud[39154]=16'h3572;
aud[39155]=16'h357e;
aud[39156]=16'h358a;
aud[39157]=16'h3595;
aud[39158]=16'h35a1;
aud[39159]=16'h35ad;
aud[39160]=16'h35b8;
aud[39161]=16'h35c4;
aud[39162]=16'h35d0;
aud[39163]=16'h35db;
aud[39164]=16'h35e7;
aud[39165]=16'h35f2;
aud[39166]=16'h35fe;
aud[39167]=16'h3609;
aud[39168]=16'h3615;
aud[39169]=16'h3620;
aud[39170]=16'h362c;
aud[39171]=16'h3637;
aud[39172]=16'h3643;
aud[39173]=16'h364e;
aud[39174]=16'h3659;
aud[39175]=16'h3665;
aud[39176]=16'h3670;
aud[39177]=16'h367b;
aud[39178]=16'h3686;
aud[39179]=16'h3692;
aud[39180]=16'h369d;
aud[39181]=16'h36a8;
aud[39182]=16'h36b3;
aud[39183]=16'h36be;
aud[39184]=16'h36c9;
aud[39185]=16'h36d4;
aud[39186]=16'h36e0;
aud[39187]=16'h36eb;
aud[39188]=16'h36f6;
aud[39189]=16'h3701;
aud[39190]=16'h370b;
aud[39191]=16'h3716;
aud[39192]=16'h3721;
aud[39193]=16'h372c;
aud[39194]=16'h3737;
aud[39195]=16'h3742;
aud[39196]=16'h374d;
aud[39197]=16'h3757;
aud[39198]=16'h3762;
aud[39199]=16'h376d;
aud[39200]=16'h3778;
aud[39201]=16'h3782;
aud[39202]=16'h378d;
aud[39203]=16'h3798;
aud[39204]=16'h37a2;
aud[39205]=16'h37ad;
aud[39206]=16'h37b7;
aud[39207]=16'h37c2;
aud[39208]=16'h37cc;
aud[39209]=16'h37d7;
aud[39210]=16'h37e1;
aud[39211]=16'h37ec;
aud[39212]=16'h37f6;
aud[39213]=16'h3801;
aud[39214]=16'h380b;
aud[39215]=16'h3815;
aud[39216]=16'h3820;
aud[39217]=16'h382a;
aud[39218]=16'h3834;
aud[39219]=16'h383f;
aud[39220]=16'h3849;
aud[39221]=16'h3853;
aud[39222]=16'h385d;
aud[39223]=16'h3867;
aud[39224]=16'h3871;
aud[39225]=16'h387b;
aud[39226]=16'h3886;
aud[39227]=16'h3890;
aud[39228]=16'h389a;
aud[39229]=16'h38a4;
aud[39230]=16'h38ae;
aud[39231]=16'h38b8;
aud[39232]=16'h38c1;
aud[39233]=16'h38cb;
aud[39234]=16'h38d5;
aud[39235]=16'h38df;
aud[39236]=16'h38e9;
aud[39237]=16'h38f3;
aud[39238]=16'h38fd;
aud[39239]=16'h3906;
aud[39240]=16'h3910;
aud[39241]=16'h391a;
aud[39242]=16'h3923;
aud[39243]=16'h392d;
aud[39244]=16'h3937;
aud[39245]=16'h3940;
aud[39246]=16'h394a;
aud[39247]=16'h3953;
aud[39248]=16'h395d;
aud[39249]=16'h3966;
aud[39250]=16'h3970;
aud[39251]=16'h3979;
aud[39252]=16'h3983;
aud[39253]=16'h398c;
aud[39254]=16'h3995;
aud[39255]=16'h399f;
aud[39256]=16'h39a8;
aud[39257]=16'h39b1;
aud[39258]=16'h39bb;
aud[39259]=16'h39c4;
aud[39260]=16'h39cd;
aud[39261]=16'h39d6;
aud[39262]=16'h39e0;
aud[39263]=16'h39e9;
aud[39264]=16'h39f2;
aud[39265]=16'h39fb;
aud[39266]=16'h3a04;
aud[39267]=16'h3a0d;
aud[39268]=16'h3a16;
aud[39269]=16'h3a1f;
aud[39270]=16'h3a28;
aud[39271]=16'h3a31;
aud[39272]=16'h3a3a;
aud[39273]=16'h3a43;
aud[39274]=16'h3a4c;
aud[39275]=16'h3a54;
aud[39276]=16'h3a5d;
aud[39277]=16'h3a66;
aud[39278]=16'h3a6f;
aud[39279]=16'h3a78;
aud[39280]=16'h3a80;
aud[39281]=16'h3a89;
aud[39282]=16'h3a92;
aud[39283]=16'h3a9a;
aud[39284]=16'h3aa3;
aud[39285]=16'h3aab;
aud[39286]=16'h3ab4;
aud[39287]=16'h3abc;
aud[39288]=16'h3ac5;
aud[39289]=16'h3acd;
aud[39290]=16'h3ad6;
aud[39291]=16'h3ade;
aud[39292]=16'h3ae7;
aud[39293]=16'h3aef;
aud[39294]=16'h3af7;
aud[39295]=16'h3b00;
aud[39296]=16'h3b08;
aud[39297]=16'h3b10;
aud[39298]=16'h3b19;
aud[39299]=16'h3b21;
aud[39300]=16'h3b29;
aud[39301]=16'h3b31;
aud[39302]=16'h3b39;
aud[39303]=16'h3b41;
aud[39304]=16'h3b4a;
aud[39305]=16'h3b52;
aud[39306]=16'h3b5a;
aud[39307]=16'h3b62;
aud[39308]=16'h3b6a;
aud[39309]=16'h3b72;
aud[39310]=16'h3b7a;
aud[39311]=16'h3b81;
aud[39312]=16'h3b89;
aud[39313]=16'h3b91;
aud[39314]=16'h3b99;
aud[39315]=16'h3ba1;
aud[39316]=16'h3ba9;
aud[39317]=16'h3bb0;
aud[39318]=16'h3bb8;
aud[39319]=16'h3bc0;
aud[39320]=16'h3bc7;
aud[39321]=16'h3bcf;
aud[39322]=16'h3bd7;
aud[39323]=16'h3bde;
aud[39324]=16'h3be6;
aud[39325]=16'h3bed;
aud[39326]=16'h3bf5;
aud[39327]=16'h3bfc;
aud[39328]=16'h3c04;
aud[39329]=16'h3c0b;
aud[39330]=16'h3c13;
aud[39331]=16'h3c1a;
aud[39332]=16'h3c21;
aud[39333]=16'h3c29;
aud[39334]=16'h3c30;
aud[39335]=16'h3c37;
aud[39336]=16'h3c3f;
aud[39337]=16'h3c46;
aud[39338]=16'h3c4d;
aud[39339]=16'h3c54;
aud[39340]=16'h3c5b;
aud[39341]=16'h3c63;
aud[39342]=16'h3c6a;
aud[39343]=16'h3c71;
aud[39344]=16'h3c78;
aud[39345]=16'h3c7f;
aud[39346]=16'h3c86;
aud[39347]=16'h3c8d;
aud[39348]=16'h3c94;
aud[39349]=16'h3c9b;
aud[39350]=16'h3ca1;
aud[39351]=16'h3ca8;
aud[39352]=16'h3caf;
aud[39353]=16'h3cb6;
aud[39354]=16'h3cbd;
aud[39355]=16'h3cc3;
aud[39356]=16'h3cca;
aud[39357]=16'h3cd1;
aud[39358]=16'h3cd7;
aud[39359]=16'h3cde;
aud[39360]=16'h3ce5;
aud[39361]=16'h3ceb;
aud[39362]=16'h3cf2;
aud[39363]=16'h3cf8;
aud[39364]=16'h3cff;
aud[39365]=16'h3d05;
aud[39366]=16'h3d0c;
aud[39367]=16'h3d12;
aud[39368]=16'h3d19;
aud[39369]=16'h3d1f;
aud[39370]=16'h3d25;
aud[39371]=16'h3d2c;
aud[39372]=16'h3d32;
aud[39373]=16'h3d38;
aud[39374]=16'h3d3f;
aud[39375]=16'h3d45;
aud[39376]=16'h3d4b;
aud[39377]=16'h3d51;
aud[39378]=16'h3d57;
aud[39379]=16'h3d5d;
aud[39380]=16'h3d63;
aud[39381]=16'h3d69;
aud[39382]=16'h3d6f;
aud[39383]=16'h3d75;
aud[39384]=16'h3d7b;
aud[39385]=16'h3d81;
aud[39386]=16'h3d87;
aud[39387]=16'h3d8d;
aud[39388]=16'h3d93;
aud[39389]=16'h3d99;
aud[39390]=16'h3d9f;
aud[39391]=16'h3da4;
aud[39392]=16'h3daa;
aud[39393]=16'h3db0;
aud[39394]=16'h3db6;
aud[39395]=16'h3dbb;
aud[39396]=16'h3dc1;
aud[39397]=16'h3dc7;
aud[39398]=16'h3dcc;
aud[39399]=16'h3dd2;
aud[39400]=16'h3dd7;
aud[39401]=16'h3ddd;
aud[39402]=16'h3de2;
aud[39403]=16'h3de8;
aud[39404]=16'h3ded;
aud[39405]=16'h3df3;
aud[39406]=16'h3df8;
aud[39407]=16'h3dfd;
aud[39408]=16'h3e03;
aud[39409]=16'h3e08;
aud[39410]=16'h3e0d;
aud[39411]=16'h3e12;
aud[39412]=16'h3e18;
aud[39413]=16'h3e1d;
aud[39414]=16'h3e22;
aud[39415]=16'h3e27;
aud[39416]=16'h3e2c;
aud[39417]=16'h3e31;
aud[39418]=16'h3e36;
aud[39419]=16'h3e3b;
aud[39420]=16'h3e40;
aud[39421]=16'h3e45;
aud[39422]=16'h3e4a;
aud[39423]=16'h3e4f;
aud[39424]=16'h3e54;
aud[39425]=16'h3e59;
aud[39426]=16'h3e5e;
aud[39427]=16'h3e62;
aud[39428]=16'h3e67;
aud[39429]=16'h3e6c;
aud[39430]=16'h3e71;
aud[39431]=16'h3e75;
aud[39432]=16'h3e7a;
aud[39433]=16'h3e7f;
aud[39434]=16'h3e83;
aud[39435]=16'h3e88;
aud[39436]=16'h3e8c;
aud[39437]=16'h3e91;
aud[39438]=16'h3e95;
aud[39439]=16'h3e9a;
aud[39440]=16'h3e9e;
aud[39441]=16'h3ea3;
aud[39442]=16'h3ea7;
aud[39443]=16'h3eac;
aud[39444]=16'h3eb0;
aud[39445]=16'h3eb4;
aud[39446]=16'h3eb9;
aud[39447]=16'h3ebd;
aud[39448]=16'h3ec1;
aud[39449]=16'h3ec5;
aud[39450]=16'h3ec9;
aud[39451]=16'h3ecd;
aud[39452]=16'h3ed2;
aud[39453]=16'h3ed6;
aud[39454]=16'h3eda;
aud[39455]=16'h3ede;
aud[39456]=16'h3ee2;
aud[39457]=16'h3ee6;
aud[39458]=16'h3eea;
aud[39459]=16'h3eee;
aud[39460]=16'h3ef2;
aud[39461]=16'h3ef5;
aud[39462]=16'h3ef9;
aud[39463]=16'h3efd;
aud[39464]=16'h3f01;
aud[39465]=16'h3f05;
aud[39466]=16'h3f08;
aud[39467]=16'h3f0c;
aud[39468]=16'h3f10;
aud[39469]=16'h3f13;
aud[39470]=16'h3f17;
aud[39471]=16'h3f1b;
aud[39472]=16'h3f1e;
aud[39473]=16'h3f22;
aud[39474]=16'h3f25;
aud[39475]=16'h3f29;
aud[39476]=16'h3f2c;
aud[39477]=16'h3f30;
aud[39478]=16'h3f33;
aud[39479]=16'h3f36;
aud[39480]=16'h3f3a;
aud[39481]=16'h3f3d;
aud[39482]=16'h3f40;
aud[39483]=16'h3f43;
aud[39484]=16'h3f47;
aud[39485]=16'h3f4a;
aud[39486]=16'h3f4d;
aud[39487]=16'h3f50;
aud[39488]=16'h3f53;
aud[39489]=16'h3f56;
aud[39490]=16'h3f5a;
aud[39491]=16'h3f5d;
aud[39492]=16'h3f60;
aud[39493]=16'h3f63;
aud[39494]=16'h3f65;
aud[39495]=16'h3f68;
aud[39496]=16'h3f6b;
aud[39497]=16'h3f6e;
aud[39498]=16'h3f71;
aud[39499]=16'h3f74;
aud[39500]=16'h3f77;
aud[39501]=16'h3f79;
aud[39502]=16'h3f7c;
aud[39503]=16'h3f7f;
aud[39504]=16'h3f81;
aud[39505]=16'h3f84;
aud[39506]=16'h3f87;
aud[39507]=16'h3f89;
aud[39508]=16'h3f8c;
aud[39509]=16'h3f8e;
aud[39510]=16'h3f91;
aud[39511]=16'h3f93;
aud[39512]=16'h3f96;
aud[39513]=16'h3f98;
aud[39514]=16'h3f9b;
aud[39515]=16'h3f9d;
aud[39516]=16'h3f9f;
aud[39517]=16'h3fa2;
aud[39518]=16'h3fa4;
aud[39519]=16'h3fa6;
aud[39520]=16'h3fa8;
aud[39521]=16'h3fab;
aud[39522]=16'h3fad;
aud[39523]=16'h3faf;
aud[39524]=16'h3fb1;
aud[39525]=16'h3fb3;
aud[39526]=16'h3fb5;
aud[39527]=16'h3fb7;
aud[39528]=16'h3fb9;
aud[39529]=16'h3fbb;
aud[39530]=16'h3fbd;
aud[39531]=16'h3fbf;
aud[39532]=16'h3fc1;
aud[39533]=16'h3fc3;
aud[39534]=16'h3fc5;
aud[39535]=16'h3fc7;
aud[39536]=16'h3fc8;
aud[39537]=16'h3fca;
aud[39538]=16'h3fcc;
aud[39539]=16'h3fcd;
aud[39540]=16'h3fcf;
aud[39541]=16'h3fd1;
aud[39542]=16'h3fd2;
aud[39543]=16'h3fd4;
aud[39544]=16'h3fd6;
aud[39545]=16'h3fd7;
aud[39546]=16'h3fd9;
aud[39547]=16'h3fda;
aud[39548]=16'h3fdc;
aud[39549]=16'h3fdd;
aud[39550]=16'h3fde;
aud[39551]=16'h3fe0;
aud[39552]=16'h3fe1;
aud[39553]=16'h3fe2;
aud[39554]=16'h3fe4;
aud[39555]=16'h3fe5;
aud[39556]=16'h3fe6;
aud[39557]=16'h3fe7;
aud[39558]=16'h3fe8;
aud[39559]=16'h3fea;
aud[39560]=16'h3feb;
aud[39561]=16'h3fec;
aud[39562]=16'h3fed;
aud[39563]=16'h3fee;
aud[39564]=16'h3fef;
aud[39565]=16'h3ff0;
aud[39566]=16'h3ff1;
aud[39567]=16'h3ff2;
aud[39568]=16'h3ff3;
aud[39569]=16'h3ff3;
aud[39570]=16'h3ff4;
aud[39571]=16'h3ff5;
aud[39572]=16'h3ff6;
aud[39573]=16'h3ff7;
aud[39574]=16'h3ff7;
aud[39575]=16'h3ff8;
aud[39576]=16'h3ff9;
aud[39577]=16'h3ff9;
aud[39578]=16'h3ffa;
aud[39579]=16'h3ffa;
aud[39580]=16'h3ffb;
aud[39581]=16'h3ffb;
aud[39582]=16'h3ffc;
aud[39583]=16'h3ffc;
aud[39584]=16'h3ffd;
aud[39585]=16'h3ffd;
aud[39586]=16'h3ffe;
aud[39587]=16'h3ffe;
aud[39588]=16'h3ffe;
aud[39589]=16'h3fff;
aud[39590]=16'h3fff;
aud[39591]=16'h3fff;
aud[39592]=16'h3fff;
aud[39593]=16'h3fff;
aud[39594]=16'h4000;
aud[39595]=16'h4000;
aud[39596]=16'h4000;
aud[39597]=16'h4000;
aud[39598]=16'h4000;
aud[39599]=16'h4000;
aud[39600]=16'h4000;
aud[39601]=16'h4000;
aud[39602]=16'h4000;
aud[39603]=16'h4000;
aud[39604]=16'h4000;
aud[39605]=16'h3fff;
aud[39606]=16'h3fff;
aud[39607]=16'h3fff;
aud[39608]=16'h3fff;
aud[39609]=16'h3fff;
aud[39610]=16'h3ffe;
aud[39611]=16'h3ffe;
aud[39612]=16'h3ffe;
aud[39613]=16'h3ffd;
aud[39614]=16'h3ffd;
aud[39615]=16'h3ffc;
aud[39616]=16'h3ffc;
aud[39617]=16'h3ffb;
aud[39618]=16'h3ffb;
aud[39619]=16'h3ffa;
aud[39620]=16'h3ffa;
aud[39621]=16'h3ff9;
aud[39622]=16'h3ff9;
aud[39623]=16'h3ff8;
aud[39624]=16'h3ff7;
aud[39625]=16'h3ff7;
aud[39626]=16'h3ff6;
aud[39627]=16'h3ff5;
aud[39628]=16'h3ff4;
aud[39629]=16'h3ff3;
aud[39630]=16'h3ff3;
aud[39631]=16'h3ff2;
aud[39632]=16'h3ff1;
aud[39633]=16'h3ff0;
aud[39634]=16'h3fef;
aud[39635]=16'h3fee;
aud[39636]=16'h3fed;
aud[39637]=16'h3fec;
aud[39638]=16'h3feb;
aud[39639]=16'h3fea;
aud[39640]=16'h3fe8;
aud[39641]=16'h3fe7;
aud[39642]=16'h3fe6;
aud[39643]=16'h3fe5;
aud[39644]=16'h3fe4;
aud[39645]=16'h3fe2;
aud[39646]=16'h3fe1;
aud[39647]=16'h3fe0;
aud[39648]=16'h3fde;
aud[39649]=16'h3fdd;
aud[39650]=16'h3fdc;
aud[39651]=16'h3fda;
aud[39652]=16'h3fd9;
aud[39653]=16'h3fd7;
aud[39654]=16'h3fd6;
aud[39655]=16'h3fd4;
aud[39656]=16'h3fd2;
aud[39657]=16'h3fd1;
aud[39658]=16'h3fcf;
aud[39659]=16'h3fcd;
aud[39660]=16'h3fcc;
aud[39661]=16'h3fca;
aud[39662]=16'h3fc8;
aud[39663]=16'h3fc7;
aud[39664]=16'h3fc5;
aud[39665]=16'h3fc3;
aud[39666]=16'h3fc1;
aud[39667]=16'h3fbf;
aud[39668]=16'h3fbd;
aud[39669]=16'h3fbb;
aud[39670]=16'h3fb9;
aud[39671]=16'h3fb7;
aud[39672]=16'h3fb5;
aud[39673]=16'h3fb3;
aud[39674]=16'h3fb1;
aud[39675]=16'h3faf;
aud[39676]=16'h3fad;
aud[39677]=16'h3fab;
aud[39678]=16'h3fa8;
aud[39679]=16'h3fa6;
aud[39680]=16'h3fa4;
aud[39681]=16'h3fa2;
aud[39682]=16'h3f9f;
aud[39683]=16'h3f9d;
aud[39684]=16'h3f9b;
aud[39685]=16'h3f98;
aud[39686]=16'h3f96;
aud[39687]=16'h3f93;
aud[39688]=16'h3f91;
aud[39689]=16'h3f8e;
aud[39690]=16'h3f8c;
aud[39691]=16'h3f89;
aud[39692]=16'h3f87;
aud[39693]=16'h3f84;
aud[39694]=16'h3f81;
aud[39695]=16'h3f7f;
aud[39696]=16'h3f7c;
aud[39697]=16'h3f79;
aud[39698]=16'h3f77;
aud[39699]=16'h3f74;
aud[39700]=16'h3f71;
aud[39701]=16'h3f6e;
aud[39702]=16'h3f6b;
aud[39703]=16'h3f68;
aud[39704]=16'h3f65;
aud[39705]=16'h3f63;
aud[39706]=16'h3f60;
aud[39707]=16'h3f5d;
aud[39708]=16'h3f5a;
aud[39709]=16'h3f56;
aud[39710]=16'h3f53;
aud[39711]=16'h3f50;
aud[39712]=16'h3f4d;
aud[39713]=16'h3f4a;
aud[39714]=16'h3f47;
aud[39715]=16'h3f43;
aud[39716]=16'h3f40;
aud[39717]=16'h3f3d;
aud[39718]=16'h3f3a;
aud[39719]=16'h3f36;
aud[39720]=16'h3f33;
aud[39721]=16'h3f30;
aud[39722]=16'h3f2c;
aud[39723]=16'h3f29;
aud[39724]=16'h3f25;
aud[39725]=16'h3f22;
aud[39726]=16'h3f1e;
aud[39727]=16'h3f1b;
aud[39728]=16'h3f17;
aud[39729]=16'h3f13;
aud[39730]=16'h3f10;
aud[39731]=16'h3f0c;
aud[39732]=16'h3f08;
aud[39733]=16'h3f05;
aud[39734]=16'h3f01;
aud[39735]=16'h3efd;
aud[39736]=16'h3ef9;
aud[39737]=16'h3ef5;
aud[39738]=16'h3ef2;
aud[39739]=16'h3eee;
aud[39740]=16'h3eea;
aud[39741]=16'h3ee6;
aud[39742]=16'h3ee2;
aud[39743]=16'h3ede;
aud[39744]=16'h3eda;
aud[39745]=16'h3ed6;
aud[39746]=16'h3ed2;
aud[39747]=16'h3ecd;
aud[39748]=16'h3ec9;
aud[39749]=16'h3ec5;
aud[39750]=16'h3ec1;
aud[39751]=16'h3ebd;
aud[39752]=16'h3eb9;
aud[39753]=16'h3eb4;
aud[39754]=16'h3eb0;
aud[39755]=16'h3eac;
aud[39756]=16'h3ea7;
aud[39757]=16'h3ea3;
aud[39758]=16'h3e9e;
aud[39759]=16'h3e9a;
aud[39760]=16'h3e95;
aud[39761]=16'h3e91;
aud[39762]=16'h3e8c;
aud[39763]=16'h3e88;
aud[39764]=16'h3e83;
aud[39765]=16'h3e7f;
aud[39766]=16'h3e7a;
aud[39767]=16'h3e75;
aud[39768]=16'h3e71;
aud[39769]=16'h3e6c;
aud[39770]=16'h3e67;
aud[39771]=16'h3e62;
aud[39772]=16'h3e5e;
aud[39773]=16'h3e59;
aud[39774]=16'h3e54;
aud[39775]=16'h3e4f;
aud[39776]=16'h3e4a;
aud[39777]=16'h3e45;
aud[39778]=16'h3e40;
aud[39779]=16'h3e3b;
aud[39780]=16'h3e36;
aud[39781]=16'h3e31;
aud[39782]=16'h3e2c;
aud[39783]=16'h3e27;
aud[39784]=16'h3e22;
aud[39785]=16'h3e1d;
aud[39786]=16'h3e18;
aud[39787]=16'h3e12;
aud[39788]=16'h3e0d;
aud[39789]=16'h3e08;
aud[39790]=16'h3e03;
aud[39791]=16'h3dfd;
aud[39792]=16'h3df8;
aud[39793]=16'h3df3;
aud[39794]=16'h3ded;
aud[39795]=16'h3de8;
aud[39796]=16'h3de2;
aud[39797]=16'h3ddd;
aud[39798]=16'h3dd7;
aud[39799]=16'h3dd2;
aud[39800]=16'h3dcc;
aud[39801]=16'h3dc7;
aud[39802]=16'h3dc1;
aud[39803]=16'h3dbb;
aud[39804]=16'h3db6;
aud[39805]=16'h3db0;
aud[39806]=16'h3daa;
aud[39807]=16'h3da4;
aud[39808]=16'h3d9f;
aud[39809]=16'h3d99;
aud[39810]=16'h3d93;
aud[39811]=16'h3d8d;
aud[39812]=16'h3d87;
aud[39813]=16'h3d81;
aud[39814]=16'h3d7b;
aud[39815]=16'h3d75;
aud[39816]=16'h3d6f;
aud[39817]=16'h3d69;
aud[39818]=16'h3d63;
aud[39819]=16'h3d5d;
aud[39820]=16'h3d57;
aud[39821]=16'h3d51;
aud[39822]=16'h3d4b;
aud[39823]=16'h3d45;
aud[39824]=16'h3d3f;
aud[39825]=16'h3d38;
aud[39826]=16'h3d32;
aud[39827]=16'h3d2c;
aud[39828]=16'h3d25;
aud[39829]=16'h3d1f;
aud[39830]=16'h3d19;
aud[39831]=16'h3d12;
aud[39832]=16'h3d0c;
aud[39833]=16'h3d05;
aud[39834]=16'h3cff;
aud[39835]=16'h3cf8;
aud[39836]=16'h3cf2;
aud[39837]=16'h3ceb;
aud[39838]=16'h3ce5;
aud[39839]=16'h3cde;
aud[39840]=16'h3cd7;
aud[39841]=16'h3cd1;
aud[39842]=16'h3cca;
aud[39843]=16'h3cc3;
aud[39844]=16'h3cbd;
aud[39845]=16'h3cb6;
aud[39846]=16'h3caf;
aud[39847]=16'h3ca8;
aud[39848]=16'h3ca1;
aud[39849]=16'h3c9b;
aud[39850]=16'h3c94;
aud[39851]=16'h3c8d;
aud[39852]=16'h3c86;
aud[39853]=16'h3c7f;
aud[39854]=16'h3c78;
aud[39855]=16'h3c71;
aud[39856]=16'h3c6a;
aud[39857]=16'h3c63;
aud[39858]=16'h3c5b;
aud[39859]=16'h3c54;
aud[39860]=16'h3c4d;
aud[39861]=16'h3c46;
aud[39862]=16'h3c3f;
aud[39863]=16'h3c37;
aud[39864]=16'h3c30;
aud[39865]=16'h3c29;
aud[39866]=16'h3c21;
aud[39867]=16'h3c1a;
aud[39868]=16'h3c13;
aud[39869]=16'h3c0b;
aud[39870]=16'h3c04;
aud[39871]=16'h3bfc;
aud[39872]=16'h3bf5;
aud[39873]=16'h3bed;
aud[39874]=16'h3be6;
aud[39875]=16'h3bde;
aud[39876]=16'h3bd7;
aud[39877]=16'h3bcf;
aud[39878]=16'h3bc7;
aud[39879]=16'h3bc0;
aud[39880]=16'h3bb8;
aud[39881]=16'h3bb0;
aud[39882]=16'h3ba9;
aud[39883]=16'h3ba1;
aud[39884]=16'h3b99;
aud[39885]=16'h3b91;
aud[39886]=16'h3b89;
aud[39887]=16'h3b81;
aud[39888]=16'h3b7a;
aud[39889]=16'h3b72;
aud[39890]=16'h3b6a;
aud[39891]=16'h3b62;
aud[39892]=16'h3b5a;
aud[39893]=16'h3b52;
aud[39894]=16'h3b4a;
aud[39895]=16'h3b41;
aud[39896]=16'h3b39;
aud[39897]=16'h3b31;
aud[39898]=16'h3b29;
aud[39899]=16'h3b21;
aud[39900]=16'h3b19;
aud[39901]=16'h3b10;
aud[39902]=16'h3b08;
aud[39903]=16'h3b00;
aud[39904]=16'h3af7;
aud[39905]=16'h3aef;
aud[39906]=16'h3ae7;
aud[39907]=16'h3ade;
aud[39908]=16'h3ad6;
aud[39909]=16'h3acd;
aud[39910]=16'h3ac5;
aud[39911]=16'h3abc;
aud[39912]=16'h3ab4;
aud[39913]=16'h3aab;
aud[39914]=16'h3aa3;
aud[39915]=16'h3a9a;
aud[39916]=16'h3a92;
aud[39917]=16'h3a89;
aud[39918]=16'h3a80;
aud[39919]=16'h3a78;
aud[39920]=16'h3a6f;
aud[39921]=16'h3a66;
aud[39922]=16'h3a5d;
aud[39923]=16'h3a54;
aud[39924]=16'h3a4c;
aud[39925]=16'h3a43;
aud[39926]=16'h3a3a;
aud[39927]=16'h3a31;
aud[39928]=16'h3a28;
aud[39929]=16'h3a1f;
aud[39930]=16'h3a16;
aud[39931]=16'h3a0d;
aud[39932]=16'h3a04;
aud[39933]=16'h39fb;
aud[39934]=16'h39f2;
aud[39935]=16'h39e9;
aud[39936]=16'h39e0;
aud[39937]=16'h39d6;
aud[39938]=16'h39cd;
aud[39939]=16'h39c4;
aud[39940]=16'h39bb;
aud[39941]=16'h39b1;
aud[39942]=16'h39a8;
aud[39943]=16'h399f;
aud[39944]=16'h3995;
aud[39945]=16'h398c;
aud[39946]=16'h3983;
aud[39947]=16'h3979;
aud[39948]=16'h3970;
aud[39949]=16'h3966;
aud[39950]=16'h395d;
aud[39951]=16'h3953;
aud[39952]=16'h394a;
aud[39953]=16'h3940;
aud[39954]=16'h3937;
aud[39955]=16'h392d;
aud[39956]=16'h3923;
aud[39957]=16'h391a;
aud[39958]=16'h3910;
aud[39959]=16'h3906;
aud[39960]=16'h38fd;
aud[39961]=16'h38f3;
aud[39962]=16'h38e9;
aud[39963]=16'h38df;
aud[39964]=16'h38d5;
aud[39965]=16'h38cb;
aud[39966]=16'h38c1;
aud[39967]=16'h38b8;
aud[39968]=16'h38ae;
aud[39969]=16'h38a4;
aud[39970]=16'h389a;
aud[39971]=16'h3890;
aud[39972]=16'h3886;
aud[39973]=16'h387b;
aud[39974]=16'h3871;
aud[39975]=16'h3867;
aud[39976]=16'h385d;
aud[39977]=16'h3853;
aud[39978]=16'h3849;
aud[39979]=16'h383f;
aud[39980]=16'h3834;
aud[39981]=16'h382a;
aud[39982]=16'h3820;
aud[39983]=16'h3815;
aud[39984]=16'h380b;
aud[39985]=16'h3801;
aud[39986]=16'h37f6;
aud[39987]=16'h37ec;
aud[39988]=16'h37e1;
aud[39989]=16'h37d7;
aud[39990]=16'h37cc;
aud[39991]=16'h37c2;
aud[39992]=16'h37b7;
aud[39993]=16'h37ad;
aud[39994]=16'h37a2;
aud[39995]=16'h3798;
aud[39996]=16'h378d;
aud[39997]=16'h3782;
aud[39998]=16'h3778;
aud[39999]=16'h376d;
aud[40000]=16'h3762;
aud[40001]=16'h3757;
aud[40002]=16'h374d;
aud[40003]=16'h3742;
aud[40004]=16'h3737;
aud[40005]=16'h372c;
aud[40006]=16'h3721;
aud[40007]=16'h3716;
aud[40008]=16'h370b;
aud[40009]=16'h3701;
aud[40010]=16'h36f6;
aud[40011]=16'h36eb;
aud[40012]=16'h36e0;
aud[40013]=16'h36d4;
aud[40014]=16'h36c9;
aud[40015]=16'h36be;
aud[40016]=16'h36b3;
aud[40017]=16'h36a8;
aud[40018]=16'h369d;
aud[40019]=16'h3692;
aud[40020]=16'h3686;
aud[40021]=16'h367b;
aud[40022]=16'h3670;
aud[40023]=16'h3665;
aud[40024]=16'h3659;
aud[40025]=16'h364e;
aud[40026]=16'h3643;
aud[40027]=16'h3637;
aud[40028]=16'h362c;
aud[40029]=16'h3620;
aud[40030]=16'h3615;
aud[40031]=16'h3609;
aud[40032]=16'h35fe;
aud[40033]=16'h35f2;
aud[40034]=16'h35e7;
aud[40035]=16'h35db;
aud[40036]=16'h35d0;
aud[40037]=16'h35c4;
aud[40038]=16'h35b8;
aud[40039]=16'h35ad;
aud[40040]=16'h35a1;
aud[40041]=16'h3595;
aud[40042]=16'h358a;
aud[40043]=16'h357e;
aud[40044]=16'h3572;
aud[40045]=16'h3566;
aud[40046]=16'h355a;
aud[40047]=16'h354f;
aud[40048]=16'h3543;
aud[40049]=16'h3537;
aud[40050]=16'h352b;
aud[40051]=16'h351f;
aud[40052]=16'h3513;
aud[40053]=16'h3507;
aud[40054]=16'h34fb;
aud[40055]=16'h34ef;
aud[40056]=16'h34e3;
aud[40057]=16'h34d7;
aud[40058]=16'h34cb;
aud[40059]=16'h34be;
aud[40060]=16'h34b2;
aud[40061]=16'h34a6;
aud[40062]=16'h349a;
aud[40063]=16'h348e;
aud[40064]=16'h3481;
aud[40065]=16'h3475;
aud[40066]=16'h3469;
aud[40067]=16'h345d;
aud[40068]=16'h3450;
aud[40069]=16'h3444;
aud[40070]=16'h3437;
aud[40071]=16'h342b;
aud[40072]=16'h341f;
aud[40073]=16'h3412;
aud[40074]=16'h3406;
aud[40075]=16'h33f9;
aud[40076]=16'h33ed;
aud[40077]=16'h33e0;
aud[40078]=16'h33d4;
aud[40079]=16'h33c7;
aud[40080]=16'h33ba;
aud[40081]=16'h33ae;
aud[40082]=16'h33a1;
aud[40083]=16'h3394;
aud[40084]=16'h3388;
aud[40085]=16'h337b;
aud[40086]=16'h336e;
aud[40087]=16'h3361;
aud[40088]=16'h3355;
aud[40089]=16'h3348;
aud[40090]=16'h333b;
aud[40091]=16'h332e;
aud[40092]=16'h3321;
aud[40093]=16'h3314;
aud[40094]=16'h3307;
aud[40095]=16'h32fa;
aud[40096]=16'h32ed;
aud[40097]=16'h32e0;
aud[40098]=16'h32d3;
aud[40099]=16'h32c6;
aud[40100]=16'h32b9;
aud[40101]=16'h32ac;
aud[40102]=16'h329f;
aud[40103]=16'h3292;
aud[40104]=16'h3285;
aud[40105]=16'h3278;
aud[40106]=16'h326a;
aud[40107]=16'h325d;
aud[40108]=16'h3250;
aud[40109]=16'h3243;
aud[40110]=16'h3235;
aud[40111]=16'h3228;
aud[40112]=16'h321b;
aud[40113]=16'h320d;
aud[40114]=16'h3200;
aud[40115]=16'h31f3;
aud[40116]=16'h31e5;
aud[40117]=16'h31d8;
aud[40118]=16'h31ca;
aud[40119]=16'h31bd;
aud[40120]=16'h31af;
aud[40121]=16'h31a2;
aud[40122]=16'h3194;
aud[40123]=16'h3187;
aud[40124]=16'h3179;
aud[40125]=16'h316b;
aud[40126]=16'h315e;
aud[40127]=16'h3150;
aud[40128]=16'h3142;
aud[40129]=16'h3135;
aud[40130]=16'h3127;
aud[40131]=16'h3119;
aud[40132]=16'h310b;
aud[40133]=16'h30fe;
aud[40134]=16'h30f0;
aud[40135]=16'h30e2;
aud[40136]=16'h30d4;
aud[40137]=16'h30c6;
aud[40138]=16'h30b8;
aud[40139]=16'h30aa;
aud[40140]=16'h309d;
aud[40141]=16'h308f;
aud[40142]=16'h3081;
aud[40143]=16'h3073;
aud[40144]=16'h3065;
aud[40145]=16'h3057;
aud[40146]=16'h3048;
aud[40147]=16'h303a;
aud[40148]=16'h302c;
aud[40149]=16'h301e;
aud[40150]=16'h3010;
aud[40151]=16'h3002;
aud[40152]=16'h2ff4;
aud[40153]=16'h2fe5;
aud[40154]=16'h2fd7;
aud[40155]=16'h2fc9;
aud[40156]=16'h2fbb;
aud[40157]=16'h2fac;
aud[40158]=16'h2f9e;
aud[40159]=16'h2f90;
aud[40160]=16'h2f81;
aud[40161]=16'h2f73;
aud[40162]=16'h2f65;
aud[40163]=16'h2f56;
aud[40164]=16'h2f48;
aud[40165]=16'h2f39;
aud[40166]=16'h2f2b;
aud[40167]=16'h2f1c;
aud[40168]=16'h2f0e;
aud[40169]=16'h2eff;
aud[40170]=16'h2ef1;
aud[40171]=16'h2ee2;
aud[40172]=16'h2ed3;
aud[40173]=16'h2ec5;
aud[40174]=16'h2eb6;
aud[40175]=16'h2ea7;
aud[40176]=16'h2e99;
aud[40177]=16'h2e8a;
aud[40178]=16'h2e7b;
aud[40179]=16'h2e6d;
aud[40180]=16'h2e5e;
aud[40181]=16'h2e4f;
aud[40182]=16'h2e40;
aud[40183]=16'h2e31;
aud[40184]=16'h2e22;
aud[40185]=16'h2e14;
aud[40186]=16'h2e05;
aud[40187]=16'h2df6;
aud[40188]=16'h2de7;
aud[40189]=16'h2dd8;
aud[40190]=16'h2dc9;
aud[40191]=16'h2dba;
aud[40192]=16'h2dab;
aud[40193]=16'h2d9c;
aud[40194]=16'h2d8d;
aud[40195]=16'h2d7e;
aud[40196]=16'h2d6f;
aud[40197]=16'h2d60;
aud[40198]=16'h2d50;
aud[40199]=16'h2d41;
aud[40200]=16'h2d32;
aud[40201]=16'h2d23;
aud[40202]=16'h2d14;
aud[40203]=16'h2d04;
aud[40204]=16'h2cf5;
aud[40205]=16'h2ce6;
aud[40206]=16'h2cd7;
aud[40207]=16'h2cc7;
aud[40208]=16'h2cb8;
aud[40209]=16'h2ca9;
aud[40210]=16'h2c99;
aud[40211]=16'h2c8a;
aud[40212]=16'h2c7a;
aud[40213]=16'h2c6b;
aud[40214]=16'h2c5c;
aud[40215]=16'h2c4c;
aud[40216]=16'h2c3d;
aud[40217]=16'h2c2d;
aud[40218]=16'h2c1e;
aud[40219]=16'h2c0e;
aud[40220]=16'h2bfe;
aud[40221]=16'h2bef;
aud[40222]=16'h2bdf;
aud[40223]=16'h2bd0;
aud[40224]=16'h2bc0;
aud[40225]=16'h2bb0;
aud[40226]=16'h2ba1;
aud[40227]=16'h2b91;
aud[40228]=16'h2b81;
aud[40229]=16'h2b71;
aud[40230]=16'h2b62;
aud[40231]=16'h2b52;
aud[40232]=16'h2b42;
aud[40233]=16'h2b32;
aud[40234]=16'h2b22;
aud[40235]=16'h2b13;
aud[40236]=16'h2b03;
aud[40237]=16'h2af3;
aud[40238]=16'h2ae3;
aud[40239]=16'h2ad3;
aud[40240]=16'h2ac3;
aud[40241]=16'h2ab3;
aud[40242]=16'h2aa3;
aud[40243]=16'h2a93;
aud[40244]=16'h2a83;
aud[40245]=16'h2a73;
aud[40246]=16'h2a63;
aud[40247]=16'h2a53;
aud[40248]=16'h2a43;
aud[40249]=16'h2a33;
aud[40250]=16'h2a23;
aud[40251]=16'h2a12;
aud[40252]=16'h2a02;
aud[40253]=16'h29f2;
aud[40254]=16'h29e2;
aud[40255]=16'h29d2;
aud[40256]=16'h29c1;
aud[40257]=16'h29b1;
aud[40258]=16'h29a1;
aud[40259]=16'h2991;
aud[40260]=16'h2980;
aud[40261]=16'h2970;
aud[40262]=16'h2960;
aud[40263]=16'h294f;
aud[40264]=16'h293f;
aud[40265]=16'h292e;
aud[40266]=16'h291e;
aud[40267]=16'h290e;
aud[40268]=16'h28fd;
aud[40269]=16'h28ed;
aud[40270]=16'h28dc;
aud[40271]=16'h28cc;
aud[40272]=16'h28bb;
aud[40273]=16'h28aa;
aud[40274]=16'h289a;
aud[40275]=16'h2889;
aud[40276]=16'h2879;
aud[40277]=16'h2868;
aud[40278]=16'h2857;
aud[40279]=16'h2847;
aud[40280]=16'h2836;
aud[40281]=16'h2825;
aud[40282]=16'h2815;
aud[40283]=16'h2804;
aud[40284]=16'h27f3;
aud[40285]=16'h27e2;
aud[40286]=16'h27d2;
aud[40287]=16'h27c1;
aud[40288]=16'h27b0;
aud[40289]=16'h279f;
aud[40290]=16'h278e;
aud[40291]=16'h277e;
aud[40292]=16'h276d;
aud[40293]=16'h275c;
aud[40294]=16'h274b;
aud[40295]=16'h273a;
aud[40296]=16'h2729;
aud[40297]=16'h2718;
aud[40298]=16'h2707;
aud[40299]=16'h26f6;
aud[40300]=16'h26e5;
aud[40301]=16'h26d4;
aud[40302]=16'h26c3;
aud[40303]=16'h26b2;
aud[40304]=16'h26a1;
aud[40305]=16'h2690;
aud[40306]=16'h267e;
aud[40307]=16'h266d;
aud[40308]=16'h265c;
aud[40309]=16'h264b;
aud[40310]=16'h263a;
aud[40311]=16'h2629;
aud[40312]=16'h2617;
aud[40313]=16'h2606;
aud[40314]=16'h25f5;
aud[40315]=16'h25e4;
aud[40316]=16'h25d2;
aud[40317]=16'h25c1;
aud[40318]=16'h25b0;
aud[40319]=16'h259e;
aud[40320]=16'h258d;
aud[40321]=16'h257c;
aud[40322]=16'h256a;
aud[40323]=16'h2559;
aud[40324]=16'h2547;
aud[40325]=16'h2536;
aud[40326]=16'h2524;
aud[40327]=16'h2513;
aud[40328]=16'h2501;
aud[40329]=16'h24f0;
aud[40330]=16'h24de;
aud[40331]=16'h24cd;
aud[40332]=16'h24bb;
aud[40333]=16'h24aa;
aud[40334]=16'h2498;
aud[40335]=16'h2487;
aud[40336]=16'h2475;
aud[40337]=16'h2463;
aud[40338]=16'h2452;
aud[40339]=16'h2440;
aud[40340]=16'h242e;
aud[40341]=16'h241d;
aud[40342]=16'h240b;
aud[40343]=16'h23f9;
aud[40344]=16'h23e7;
aud[40345]=16'h23d6;
aud[40346]=16'h23c4;
aud[40347]=16'h23b2;
aud[40348]=16'h23a0;
aud[40349]=16'h238e;
aud[40350]=16'h237d;
aud[40351]=16'h236b;
aud[40352]=16'h2359;
aud[40353]=16'h2347;
aud[40354]=16'h2335;
aud[40355]=16'h2323;
aud[40356]=16'h2311;
aud[40357]=16'h22ff;
aud[40358]=16'h22ed;
aud[40359]=16'h22db;
aud[40360]=16'h22c9;
aud[40361]=16'h22b7;
aud[40362]=16'h22a5;
aud[40363]=16'h2293;
aud[40364]=16'h2281;
aud[40365]=16'h226f;
aud[40366]=16'h225d;
aud[40367]=16'h224b;
aud[40368]=16'h2239;
aud[40369]=16'h2227;
aud[40370]=16'h2215;
aud[40371]=16'h2202;
aud[40372]=16'h21f0;
aud[40373]=16'h21de;
aud[40374]=16'h21cc;
aud[40375]=16'h21ba;
aud[40376]=16'h21a7;
aud[40377]=16'h2195;
aud[40378]=16'h2183;
aud[40379]=16'h2171;
aud[40380]=16'h215e;
aud[40381]=16'h214c;
aud[40382]=16'h213a;
aud[40383]=16'h2127;
aud[40384]=16'h2115;
aud[40385]=16'h2103;
aud[40386]=16'h20f0;
aud[40387]=16'h20de;
aud[40388]=16'h20cb;
aud[40389]=16'h20b9;
aud[40390]=16'h20a7;
aud[40391]=16'h2094;
aud[40392]=16'h2082;
aud[40393]=16'h206f;
aud[40394]=16'h205d;
aud[40395]=16'h204a;
aud[40396]=16'h2038;
aud[40397]=16'h2025;
aud[40398]=16'h2013;
aud[40399]=16'h2000;
aud[40400]=16'h1fed;
aud[40401]=16'h1fdb;
aud[40402]=16'h1fc8;
aud[40403]=16'h1fb6;
aud[40404]=16'h1fa3;
aud[40405]=16'h1f90;
aud[40406]=16'h1f7e;
aud[40407]=16'h1f6b;
aud[40408]=16'h1f58;
aud[40409]=16'h1f46;
aud[40410]=16'h1f33;
aud[40411]=16'h1f20;
aud[40412]=16'h1f0d;
aud[40413]=16'h1efb;
aud[40414]=16'h1ee8;
aud[40415]=16'h1ed5;
aud[40416]=16'h1ec2;
aud[40417]=16'h1eaf;
aud[40418]=16'h1e9d;
aud[40419]=16'h1e8a;
aud[40420]=16'h1e77;
aud[40421]=16'h1e64;
aud[40422]=16'h1e51;
aud[40423]=16'h1e3e;
aud[40424]=16'h1e2b;
aud[40425]=16'h1e18;
aud[40426]=16'h1e06;
aud[40427]=16'h1df3;
aud[40428]=16'h1de0;
aud[40429]=16'h1dcd;
aud[40430]=16'h1dba;
aud[40431]=16'h1da7;
aud[40432]=16'h1d94;
aud[40433]=16'h1d81;
aud[40434]=16'h1d6e;
aud[40435]=16'h1d5b;
aud[40436]=16'h1d47;
aud[40437]=16'h1d34;
aud[40438]=16'h1d21;
aud[40439]=16'h1d0e;
aud[40440]=16'h1cfb;
aud[40441]=16'h1ce8;
aud[40442]=16'h1cd5;
aud[40443]=16'h1cc2;
aud[40444]=16'h1cae;
aud[40445]=16'h1c9b;
aud[40446]=16'h1c88;
aud[40447]=16'h1c75;
aud[40448]=16'h1c62;
aud[40449]=16'h1c4e;
aud[40450]=16'h1c3b;
aud[40451]=16'h1c28;
aud[40452]=16'h1c15;
aud[40453]=16'h1c01;
aud[40454]=16'h1bee;
aud[40455]=16'h1bdb;
aud[40456]=16'h1bc8;
aud[40457]=16'h1bb4;
aud[40458]=16'h1ba1;
aud[40459]=16'h1b8d;
aud[40460]=16'h1b7a;
aud[40461]=16'h1b67;
aud[40462]=16'h1b53;
aud[40463]=16'h1b40;
aud[40464]=16'h1b2d;
aud[40465]=16'h1b19;
aud[40466]=16'h1b06;
aud[40467]=16'h1af2;
aud[40468]=16'h1adf;
aud[40469]=16'h1acb;
aud[40470]=16'h1ab8;
aud[40471]=16'h1aa4;
aud[40472]=16'h1a91;
aud[40473]=16'h1a7d;
aud[40474]=16'h1a6a;
aud[40475]=16'h1a56;
aud[40476]=16'h1a43;
aud[40477]=16'h1a2f;
aud[40478]=16'h1a1c;
aud[40479]=16'h1a08;
aud[40480]=16'h19f4;
aud[40481]=16'h19e1;
aud[40482]=16'h19cd;
aud[40483]=16'h19ba;
aud[40484]=16'h19a6;
aud[40485]=16'h1992;
aud[40486]=16'h197f;
aud[40487]=16'h196b;
aud[40488]=16'h1957;
aud[40489]=16'h1943;
aud[40490]=16'h1930;
aud[40491]=16'h191c;
aud[40492]=16'h1908;
aud[40493]=16'h18f5;
aud[40494]=16'h18e1;
aud[40495]=16'h18cd;
aud[40496]=16'h18b9;
aud[40497]=16'h18a5;
aud[40498]=16'h1892;
aud[40499]=16'h187e;
aud[40500]=16'h186a;
aud[40501]=16'h1856;
aud[40502]=16'h1842;
aud[40503]=16'h182f;
aud[40504]=16'h181b;
aud[40505]=16'h1807;
aud[40506]=16'h17f3;
aud[40507]=16'h17df;
aud[40508]=16'h17cb;
aud[40509]=16'h17b7;
aud[40510]=16'h17a3;
aud[40511]=16'h178f;
aud[40512]=16'h177b;
aud[40513]=16'h1767;
aud[40514]=16'h1753;
aud[40515]=16'h1740;
aud[40516]=16'h172c;
aud[40517]=16'h1718;
aud[40518]=16'h1704;
aud[40519]=16'h16f0;
aud[40520]=16'h16db;
aud[40521]=16'h16c7;
aud[40522]=16'h16b3;
aud[40523]=16'h169f;
aud[40524]=16'h168b;
aud[40525]=16'h1677;
aud[40526]=16'h1663;
aud[40527]=16'h164f;
aud[40528]=16'h163b;
aud[40529]=16'h1627;
aud[40530]=16'h1613;
aud[40531]=16'h15ff;
aud[40532]=16'h15ea;
aud[40533]=16'h15d6;
aud[40534]=16'h15c2;
aud[40535]=16'h15ae;
aud[40536]=16'h159a;
aud[40537]=16'h1586;
aud[40538]=16'h1571;
aud[40539]=16'h155d;
aud[40540]=16'h1549;
aud[40541]=16'h1535;
aud[40542]=16'h1520;
aud[40543]=16'h150c;
aud[40544]=16'h14f8;
aud[40545]=16'h14e4;
aud[40546]=16'h14cf;
aud[40547]=16'h14bb;
aud[40548]=16'h14a7;
aud[40549]=16'h1492;
aud[40550]=16'h147e;
aud[40551]=16'h146a;
aud[40552]=16'h1455;
aud[40553]=16'h1441;
aud[40554]=16'h142d;
aud[40555]=16'h1418;
aud[40556]=16'h1404;
aud[40557]=16'h13f0;
aud[40558]=16'h13db;
aud[40559]=16'h13c7;
aud[40560]=16'h13b3;
aud[40561]=16'h139e;
aud[40562]=16'h138a;
aud[40563]=16'h1375;
aud[40564]=16'h1361;
aud[40565]=16'h134c;
aud[40566]=16'h1338;
aud[40567]=16'h1323;
aud[40568]=16'h130f;
aud[40569]=16'h12fb;
aud[40570]=16'h12e6;
aud[40571]=16'h12d2;
aud[40572]=16'h12bd;
aud[40573]=16'h12a9;
aud[40574]=16'h1294;
aud[40575]=16'h127f;
aud[40576]=16'h126b;
aud[40577]=16'h1256;
aud[40578]=16'h1242;
aud[40579]=16'h122d;
aud[40580]=16'h1219;
aud[40581]=16'h1204;
aud[40582]=16'h11f0;
aud[40583]=16'h11db;
aud[40584]=16'h11c6;
aud[40585]=16'h11b2;
aud[40586]=16'h119d;
aud[40587]=16'h1189;
aud[40588]=16'h1174;
aud[40589]=16'h115f;
aud[40590]=16'h114b;
aud[40591]=16'h1136;
aud[40592]=16'h1121;
aud[40593]=16'h110d;
aud[40594]=16'h10f8;
aud[40595]=16'h10e3;
aud[40596]=16'h10cf;
aud[40597]=16'h10ba;
aud[40598]=16'h10a5;
aud[40599]=16'h1090;
aud[40600]=16'h107c;
aud[40601]=16'h1067;
aud[40602]=16'h1052;
aud[40603]=16'h103e;
aud[40604]=16'h1029;
aud[40605]=16'h1014;
aud[40606]=16'hfff;
aud[40607]=16'hfeb;
aud[40608]=16'hfd6;
aud[40609]=16'hfc1;
aud[40610]=16'hfac;
aud[40611]=16'hf97;
aud[40612]=16'hf83;
aud[40613]=16'hf6e;
aud[40614]=16'hf59;
aud[40615]=16'hf44;
aud[40616]=16'hf2f;
aud[40617]=16'hf1a;
aud[40618]=16'hf06;
aud[40619]=16'hef1;
aud[40620]=16'hedc;
aud[40621]=16'hec7;
aud[40622]=16'heb2;
aud[40623]=16'he9d;
aud[40624]=16'he88;
aud[40625]=16'he74;
aud[40626]=16'he5f;
aud[40627]=16'he4a;
aud[40628]=16'he35;
aud[40629]=16'he20;
aud[40630]=16'he0b;
aud[40631]=16'hdf6;
aud[40632]=16'hde1;
aud[40633]=16'hdcc;
aud[40634]=16'hdb7;
aud[40635]=16'hda2;
aud[40636]=16'hd8d;
aud[40637]=16'hd78;
aud[40638]=16'hd63;
aud[40639]=16'hd4e;
aud[40640]=16'hd39;
aud[40641]=16'hd24;
aud[40642]=16'hd0f;
aud[40643]=16'hcfa;
aud[40644]=16'hce5;
aud[40645]=16'hcd0;
aud[40646]=16'hcbb;
aud[40647]=16'hca6;
aud[40648]=16'hc91;
aud[40649]=16'hc7c;
aud[40650]=16'hc67;
aud[40651]=16'hc52;
aud[40652]=16'hc3d;
aud[40653]=16'hc28;
aud[40654]=16'hc13;
aud[40655]=16'hbfe;
aud[40656]=16'hbe9;
aud[40657]=16'hbd4;
aud[40658]=16'hbbf;
aud[40659]=16'hbaa;
aud[40660]=16'hb95;
aud[40661]=16'hb80;
aud[40662]=16'hb6a;
aud[40663]=16'hb55;
aud[40664]=16'hb40;
aud[40665]=16'hb2b;
aud[40666]=16'hb16;
aud[40667]=16'hb01;
aud[40668]=16'haec;
aud[40669]=16'had7;
aud[40670]=16'hac1;
aud[40671]=16'haac;
aud[40672]=16'ha97;
aud[40673]=16'ha82;
aud[40674]=16'ha6d;
aud[40675]=16'ha58;
aud[40676]=16'ha43;
aud[40677]=16'ha2d;
aud[40678]=16'ha18;
aud[40679]=16'ha03;
aud[40680]=16'h9ee;
aud[40681]=16'h9d9;
aud[40682]=16'h9c3;
aud[40683]=16'h9ae;
aud[40684]=16'h999;
aud[40685]=16'h984;
aud[40686]=16'h96f;
aud[40687]=16'h959;
aud[40688]=16'h944;
aud[40689]=16'h92f;
aud[40690]=16'h91a;
aud[40691]=16'h905;
aud[40692]=16'h8ef;
aud[40693]=16'h8da;
aud[40694]=16'h8c5;
aud[40695]=16'h8b0;
aud[40696]=16'h89a;
aud[40697]=16'h885;
aud[40698]=16'h870;
aud[40699]=16'h85b;
aud[40700]=16'h845;
aud[40701]=16'h830;
aud[40702]=16'h81b;
aud[40703]=16'h805;
aud[40704]=16'h7f0;
aud[40705]=16'h7db;
aud[40706]=16'h7c6;
aud[40707]=16'h7b0;
aud[40708]=16'h79b;
aud[40709]=16'h786;
aud[40710]=16'h770;
aud[40711]=16'h75b;
aud[40712]=16'h746;
aud[40713]=16'h731;
aud[40714]=16'h71b;
aud[40715]=16'h706;
aud[40716]=16'h6f1;
aud[40717]=16'h6db;
aud[40718]=16'h6c6;
aud[40719]=16'h6b1;
aud[40720]=16'h69b;
aud[40721]=16'h686;
aud[40722]=16'h671;
aud[40723]=16'h65b;
aud[40724]=16'h646;
aud[40725]=16'h631;
aud[40726]=16'h61b;
aud[40727]=16'h606;
aud[40728]=16'h5f1;
aud[40729]=16'h5db;
aud[40730]=16'h5c6;
aud[40731]=16'h5b0;
aud[40732]=16'h59b;
aud[40733]=16'h586;
aud[40734]=16'h570;
aud[40735]=16'h55b;
aud[40736]=16'h546;
aud[40737]=16'h530;
aud[40738]=16'h51b;
aud[40739]=16'h505;
aud[40740]=16'h4f0;
aud[40741]=16'h4db;
aud[40742]=16'h4c5;
aud[40743]=16'h4b0;
aud[40744]=16'h49b;
aud[40745]=16'h485;
aud[40746]=16'h470;
aud[40747]=16'h45a;
aud[40748]=16'h445;
aud[40749]=16'h430;
aud[40750]=16'h41a;
aud[40751]=16'h405;
aud[40752]=16'h3ef;
aud[40753]=16'h3da;
aud[40754]=16'h3c5;
aud[40755]=16'h3af;
aud[40756]=16'h39a;
aud[40757]=16'h384;
aud[40758]=16'h36f;
aud[40759]=16'h359;
aud[40760]=16'h344;
aud[40761]=16'h32f;
aud[40762]=16'h319;
aud[40763]=16'h304;
aud[40764]=16'h2ee;
aud[40765]=16'h2d9;
aud[40766]=16'h2c4;
aud[40767]=16'h2ae;
aud[40768]=16'h299;
aud[40769]=16'h283;
aud[40770]=16'h26e;
aud[40771]=16'h258;
aud[40772]=16'h243;
aud[40773]=16'h22e;
aud[40774]=16'h218;
aud[40775]=16'h203;
aud[40776]=16'h1ed;
aud[40777]=16'h1d8;
aud[40778]=16'h1c2;
aud[40779]=16'h1ad;
aud[40780]=16'h197;
aud[40781]=16'h182;
aud[40782]=16'h16d;
aud[40783]=16'h157;
aud[40784]=16'h142;
aud[40785]=16'h12c;
aud[40786]=16'h117;
aud[40787]=16'h101;
aud[40788]=16'hec;
aud[40789]=16'hd6;
aud[40790]=16'hc1;
aud[40791]=16'hac;
aud[40792]=16'h96;
aud[40793]=16'h81;
aud[40794]=16'h6b;
aud[40795]=16'h56;
aud[40796]=16'h40;
aud[40797]=16'h2b;
aud[40798]=16'h15;
aud[40799]=16'h0;
aud[40800]=16'hffeb;
aud[40801]=16'hffd5;
aud[40802]=16'hffc0;
aud[40803]=16'hffaa;
aud[40804]=16'hff95;
aud[40805]=16'hff7f;
aud[40806]=16'hff6a;
aud[40807]=16'hff54;
aud[40808]=16'hff3f;
aud[40809]=16'hff2a;
aud[40810]=16'hff14;
aud[40811]=16'hfeff;
aud[40812]=16'hfee9;
aud[40813]=16'hfed4;
aud[40814]=16'hfebe;
aud[40815]=16'hfea9;
aud[40816]=16'hfe93;
aud[40817]=16'hfe7e;
aud[40818]=16'hfe69;
aud[40819]=16'hfe53;
aud[40820]=16'hfe3e;
aud[40821]=16'hfe28;
aud[40822]=16'hfe13;
aud[40823]=16'hfdfd;
aud[40824]=16'hfde8;
aud[40825]=16'hfdd2;
aud[40826]=16'hfdbd;
aud[40827]=16'hfda8;
aud[40828]=16'hfd92;
aud[40829]=16'hfd7d;
aud[40830]=16'hfd67;
aud[40831]=16'hfd52;
aud[40832]=16'hfd3c;
aud[40833]=16'hfd27;
aud[40834]=16'hfd12;
aud[40835]=16'hfcfc;
aud[40836]=16'hfce7;
aud[40837]=16'hfcd1;
aud[40838]=16'hfcbc;
aud[40839]=16'hfca7;
aud[40840]=16'hfc91;
aud[40841]=16'hfc7c;
aud[40842]=16'hfc66;
aud[40843]=16'hfc51;
aud[40844]=16'hfc3b;
aud[40845]=16'hfc26;
aud[40846]=16'hfc11;
aud[40847]=16'hfbfb;
aud[40848]=16'hfbe6;
aud[40849]=16'hfbd0;
aud[40850]=16'hfbbb;
aud[40851]=16'hfba6;
aud[40852]=16'hfb90;
aud[40853]=16'hfb7b;
aud[40854]=16'hfb65;
aud[40855]=16'hfb50;
aud[40856]=16'hfb3b;
aud[40857]=16'hfb25;
aud[40858]=16'hfb10;
aud[40859]=16'hfafb;
aud[40860]=16'hfae5;
aud[40861]=16'hfad0;
aud[40862]=16'hfaba;
aud[40863]=16'hfaa5;
aud[40864]=16'hfa90;
aud[40865]=16'hfa7a;
aud[40866]=16'hfa65;
aud[40867]=16'hfa50;
aud[40868]=16'hfa3a;
aud[40869]=16'hfa25;
aud[40870]=16'hfa0f;
aud[40871]=16'hf9fa;
aud[40872]=16'hf9e5;
aud[40873]=16'hf9cf;
aud[40874]=16'hf9ba;
aud[40875]=16'hf9a5;
aud[40876]=16'hf98f;
aud[40877]=16'hf97a;
aud[40878]=16'hf965;
aud[40879]=16'hf94f;
aud[40880]=16'hf93a;
aud[40881]=16'hf925;
aud[40882]=16'hf90f;
aud[40883]=16'hf8fa;
aud[40884]=16'hf8e5;
aud[40885]=16'hf8cf;
aud[40886]=16'hf8ba;
aud[40887]=16'hf8a5;
aud[40888]=16'hf890;
aud[40889]=16'hf87a;
aud[40890]=16'hf865;
aud[40891]=16'hf850;
aud[40892]=16'hf83a;
aud[40893]=16'hf825;
aud[40894]=16'hf810;
aud[40895]=16'hf7fb;
aud[40896]=16'hf7e5;
aud[40897]=16'hf7d0;
aud[40898]=16'hf7bb;
aud[40899]=16'hf7a5;
aud[40900]=16'hf790;
aud[40901]=16'hf77b;
aud[40902]=16'hf766;
aud[40903]=16'hf750;
aud[40904]=16'hf73b;
aud[40905]=16'hf726;
aud[40906]=16'hf711;
aud[40907]=16'hf6fb;
aud[40908]=16'hf6e6;
aud[40909]=16'hf6d1;
aud[40910]=16'hf6bc;
aud[40911]=16'hf6a7;
aud[40912]=16'hf691;
aud[40913]=16'hf67c;
aud[40914]=16'hf667;
aud[40915]=16'hf652;
aud[40916]=16'hf63d;
aud[40917]=16'hf627;
aud[40918]=16'hf612;
aud[40919]=16'hf5fd;
aud[40920]=16'hf5e8;
aud[40921]=16'hf5d3;
aud[40922]=16'hf5bd;
aud[40923]=16'hf5a8;
aud[40924]=16'hf593;
aud[40925]=16'hf57e;
aud[40926]=16'hf569;
aud[40927]=16'hf554;
aud[40928]=16'hf53f;
aud[40929]=16'hf529;
aud[40930]=16'hf514;
aud[40931]=16'hf4ff;
aud[40932]=16'hf4ea;
aud[40933]=16'hf4d5;
aud[40934]=16'hf4c0;
aud[40935]=16'hf4ab;
aud[40936]=16'hf496;
aud[40937]=16'hf480;
aud[40938]=16'hf46b;
aud[40939]=16'hf456;
aud[40940]=16'hf441;
aud[40941]=16'hf42c;
aud[40942]=16'hf417;
aud[40943]=16'hf402;
aud[40944]=16'hf3ed;
aud[40945]=16'hf3d8;
aud[40946]=16'hf3c3;
aud[40947]=16'hf3ae;
aud[40948]=16'hf399;
aud[40949]=16'hf384;
aud[40950]=16'hf36f;
aud[40951]=16'hf35a;
aud[40952]=16'hf345;
aud[40953]=16'hf330;
aud[40954]=16'hf31b;
aud[40955]=16'hf306;
aud[40956]=16'hf2f1;
aud[40957]=16'hf2dc;
aud[40958]=16'hf2c7;
aud[40959]=16'hf2b2;
aud[40960]=16'hf29d;
aud[40961]=16'hf288;
aud[40962]=16'hf273;
aud[40963]=16'hf25e;
aud[40964]=16'hf249;
aud[40965]=16'hf234;
aud[40966]=16'hf21f;
aud[40967]=16'hf20a;
aud[40968]=16'hf1f5;
aud[40969]=16'hf1e0;
aud[40970]=16'hf1cb;
aud[40971]=16'hf1b6;
aud[40972]=16'hf1a1;
aud[40973]=16'hf18c;
aud[40974]=16'hf178;
aud[40975]=16'hf163;
aud[40976]=16'hf14e;
aud[40977]=16'hf139;
aud[40978]=16'hf124;
aud[40979]=16'hf10f;
aud[40980]=16'hf0fa;
aud[40981]=16'hf0e6;
aud[40982]=16'hf0d1;
aud[40983]=16'hf0bc;
aud[40984]=16'hf0a7;
aud[40985]=16'hf092;
aud[40986]=16'hf07d;
aud[40987]=16'hf069;
aud[40988]=16'hf054;
aud[40989]=16'hf03f;
aud[40990]=16'hf02a;
aud[40991]=16'hf015;
aud[40992]=16'hf001;
aud[40993]=16'hefec;
aud[40994]=16'hefd7;
aud[40995]=16'hefc2;
aud[40996]=16'hefae;
aud[40997]=16'hef99;
aud[40998]=16'hef84;
aud[40999]=16'hef70;
aud[41000]=16'hef5b;
aud[41001]=16'hef46;
aud[41002]=16'hef31;
aud[41003]=16'hef1d;
aud[41004]=16'hef08;
aud[41005]=16'heef3;
aud[41006]=16'heedf;
aud[41007]=16'heeca;
aud[41008]=16'heeb5;
aud[41009]=16'heea1;
aud[41010]=16'hee8c;
aud[41011]=16'hee77;
aud[41012]=16'hee63;
aud[41013]=16'hee4e;
aud[41014]=16'hee3a;
aud[41015]=16'hee25;
aud[41016]=16'hee10;
aud[41017]=16'hedfc;
aud[41018]=16'hede7;
aud[41019]=16'hedd3;
aud[41020]=16'hedbe;
aud[41021]=16'hedaa;
aud[41022]=16'hed95;
aud[41023]=16'hed81;
aud[41024]=16'hed6c;
aud[41025]=16'hed57;
aud[41026]=16'hed43;
aud[41027]=16'hed2e;
aud[41028]=16'hed1a;
aud[41029]=16'hed05;
aud[41030]=16'hecf1;
aud[41031]=16'hecdd;
aud[41032]=16'hecc8;
aud[41033]=16'hecb4;
aud[41034]=16'hec9f;
aud[41035]=16'hec8b;
aud[41036]=16'hec76;
aud[41037]=16'hec62;
aud[41038]=16'hec4d;
aud[41039]=16'hec39;
aud[41040]=16'hec25;
aud[41041]=16'hec10;
aud[41042]=16'hebfc;
aud[41043]=16'hebe8;
aud[41044]=16'hebd3;
aud[41045]=16'hebbf;
aud[41046]=16'hebab;
aud[41047]=16'heb96;
aud[41048]=16'heb82;
aud[41049]=16'heb6e;
aud[41050]=16'heb59;
aud[41051]=16'heb45;
aud[41052]=16'heb31;
aud[41053]=16'heb1c;
aud[41054]=16'heb08;
aud[41055]=16'heaf4;
aud[41056]=16'heae0;
aud[41057]=16'heacb;
aud[41058]=16'heab7;
aud[41059]=16'heaa3;
aud[41060]=16'hea8f;
aud[41061]=16'hea7a;
aud[41062]=16'hea66;
aud[41063]=16'hea52;
aud[41064]=16'hea3e;
aud[41065]=16'hea2a;
aud[41066]=16'hea16;
aud[41067]=16'hea01;
aud[41068]=16'he9ed;
aud[41069]=16'he9d9;
aud[41070]=16'he9c5;
aud[41071]=16'he9b1;
aud[41072]=16'he99d;
aud[41073]=16'he989;
aud[41074]=16'he975;
aud[41075]=16'he961;
aud[41076]=16'he94d;
aud[41077]=16'he939;
aud[41078]=16'he925;
aud[41079]=16'he910;
aud[41080]=16'he8fc;
aud[41081]=16'he8e8;
aud[41082]=16'he8d4;
aud[41083]=16'he8c0;
aud[41084]=16'he8ad;
aud[41085]=16'he899;
aud[41086]=16'he885;
aud[41087]=16'he871;
aud[41088]=16'he85d;
aud[41089]=16'he849;
aud[41090]=16'he835;
aud[41091]=16'he821;
aud[41092]=16'he80d;
aud[41093]=16'he7f9;
aud[41094]=16'he7e5;
aud[41095]=16'he7d1;
aud[41096]=16'he7be;
aud[41097]=16'he7aa;
aud[41098]=16'he796;
aud[41099]=16'he782;
aud[41100]=16'he76e;
aud[41101]=16'he75b;
aud[41102]=16'he747;
aud[41103]=16'he733;
aud[41104]=16'he71f;
aud[41105]=16'he70b;
aud[41106]=16'he6f8;
aud[41107]=16'he6e4;
aud[41108]=16'he6d0;
aud[41109]=16'he6bd;
aud[41110]=16'he6a9;
aud[41111]=16'he695;
aud[41112]=16'he681;
aud[41113]=16'he66e;
aud[41114]=16'he65a;
aud[41115]=16'he646;
aud[41116]=16'he633;
aud[41117]=16'he61f;
aud[41118]=16'he60c;
aud[41119]=16'he5f8;
aud[41120]=16'he5e4;
aud[41121]=16'he5d1;
aud[41122]=16'he5bd;
aud[41123]=16'he5aa;
aud[41124]=16'he596;
aud[41125]=16'he583;
aud[41126]=16'he56f;
aud[41127]=16'he55c;
aud[41128]=16'he548;
aud[41129]=16'he535;
aud[41130]=16'he521;
aud[41131]=16'he50e;
aud[41132]=16'he4fa;
aud[41133]=16'he4e7;
aud[41134]=16'he4d3;
aud[41135]=16'he4c0;
aud[41136]=16'he4ad;
aud[41137]=16'he499;
aud[41138]=16'he486;
aud[41139]=16'he473;
aud[41140]=16'he45f;
aud[41141]=16'he44c;
aud[41142]=16'he438;
aud[41143]=16'he425;
aud[41144]=16'he412;
aud[41145]=16'he3ff;
aud[41146]=16'he3eb;
aud[41147]=16'he3d8;
aud[41148]=16'he3c5;
aud[41149]=16'he3b2;
aud[41150]=16'he39e;
aud[41151]=16'he38b;
aud[41152]=16'he378;
aud[41153]=16'he365;
aud[41154]=16'he352;
aud[41155]=16'he33e;
aud[41156]=16'he32b;
aud[41157]=16'he318;
aud[41158]=16'he305;
aud[41159]=16'he2f2;
aud[41160]=16'he2df;
aud[41161]=16'he2cc;
aud[41162]=16'he2b9;
aud[41163]=16'he2a5;
aud[41164]=16'he292;
aud[41165]=16'he27f;
aud[41166]=16'he26c;
aud[41167]=16'he259;
aud[41168]=16'he246;
aud[41169]=16'he233;
aud[41170]=16'he220;
aud[41171]=16'he20d;
aud[41172]=16'he1fa;
aud[41173]=16'he1e8;
aud[41174]=16'he1d5;
aud[41175]=16'he1c2;
aud[41176]=16'he1af;
aud[41177]=16'he19c;
aud[41178]=16'he189;
aud[41179]=16'he176;
aud[41180]=16'he163;
aud[41181]=16'he151;
aud[41182]=16'he13e;
aud[41183]=16'he12b;
aud[41184]=16'he118;
aud[41185]=16'he105;
aud[41186]=16'he0f3;
aud[41187]=16'he0e0;
aud[41188]=16'he0cd;
aud[41189]=16'he0ba;
aud[41190]=16'he0a8;
aud[41191]=16'he095;
aud[41192]=16'he082;
aud[41193]=16'he070;
aud[41194]=16'he05d;
aud[41195]=16'he04a;
aud[41196]=16'he038;
aud[41197]=16'he025;
aud[41198]=16'he013;
aud[41199]=16'he000;
aud[41200]=16'hdfed;
aud[41201]=16'hdfdb;
aud[41202]=16'hdfc8;
aud[41203]=16'hdfb6;
aud[41204]=16'hdfa3;
aud[41205]=16'hdf91;
aud[41206]=16'hdf7e;
aud[41207]=16'hdf6c;
aud[41208]=16'hdf59;
aud[41209]=16'hdf47;
aud[41210]=16'hdf35;
aud[41211]=16'hdf22;
aud[41212]=16'hdf10;
aud[41213]=16'hdefd;
aud[41214]=16'hdeeb;
aud[41215]=16'hded9;
aud[41216]=16'hdec6;
aud[41217]=16'hdeb4;
aud[41218]=16'hdea2;
aud[41219]=16'hde8f;
aud[41220]=16'hde7d;
aud[41221]=16'hde6b;
aud[41222]=16'hde59;
aud[41223]=16'hde46;
aud[41224]=16'hde34;
aud[41225]=16'hde22;
aud[41226]=16'hde10;
aud[41227]=16'hddfe;
aud[41228]=16'hddeb;
aud[41229]=16'hddd9;
aud[41230]=16'hddc7;
aud[41231]=16'hddb5;
aud[41232]=16'hdda3;
aud[41233]=16'hdd91;
aud[41234]=16'hdd7f;
aud[41235]=16'hdd6d;
aud[41236]=16'hdd5b;
aud[41237]=16'hdd49;
aud[41238]=16'hdd37;
aud[41239]=16'hdd25;
aud[41240]=16'hdd13;
aud[41241]=16'hdd01;
aud[41242]=16'hdcef;
aud[41243]=16'hdcdd;
aud[41244]=16'hdccb;
aud[41245]=16'hdcb9;
aud[41246]=16'hdca7;
aud[41247]=16'hdc95;
aud[41248]=16'hdc83;
aud[41249]=16'hdc72;
aud[41250]=16'hdc60;
aud[41251]=16'hdc4e;
aud[41252]=16'hdc3c;
aud[41253]=16'hdc2a;
aud[41254]=16'hdc19;
aud[41255]=16'hdc07;
aud[41256]=16'hdbf5;
aud[41257]=16'hdbe3;
aud[41258]=16'hdbd2;
aud[41259]=16'hdbc0;
aud[41260]=16'hdbae;
aud[41261]=16'hdb9d;
aud[41262]=16'hdb8b;
aud[41263]=16'hdb79;
aud[41264]=16'hdb68;
aud[41265]=16'hdb56;
aud[41266]=16'hdb45;
aud[41267]=16'hdb33;
aud[41268]=16'hdb22;
aud[41269]=16'hdb10;
aud[41270]=16'hdaff;
aud[41271]=16'hdaed;
aud[41272]=16'hdadc;
aud[41273]=16'hdaca;
aud[41274]=16'hdab9;
aud[41275]=16'hdaa7;
aud[41276]=16'hda96;
aud[41277]=16'hda84;
aud[41278]=16'hda73;
aud[41279]=16'hda62;
aud[41280]=16'hda50;
aud[41281]=16'hda3f;
aud[41282]=16'hda2e;
aud[41283]=16'hda1c;
aud[41284]=16'hda0b;
aud[41285]=16'hd9fa;
aud[41286]=16'hd9e9;
aud[41287]=16'hd9d7;
aud[41288]=16'hd9c6;
aud[41289]=16'hd9b5;
aud[41290]=16'hd9a4;
aud[41291]=16'hd993;
aud[41292]=16'hd982;
aud[41293]=16'hd970;
aud[41294]=16'hd95f;
aud[41295]=16'hd94e;
aud[41296]=16'hd93d;
aud[41297]=16'hd92c;
aud[41298]=16'hd91b;
aud[41299]=16'hd90a;
aud[41300]=16'hd8f9;
aud[41301]=16'hd8e8;
aud[41302]=16'hd8d7;
aud[41303]=16'hd8c6;
aud[41304]=16'hd8b5;
aud[41305]=16'hd8a4;
aud[41306]=16'hd893;
aud[41307]=16'hd882;
aud[41308]=16'hd872;
aud[41309]=16'hd861;
aud[41310]=16'hd850;
aud[41311]=16'hd83f;
aud[41312]=16'hd82e;
aud[41313]=16'hd81e;
aud[41314]=16'hd80d;
aud[41315]=16'hd7fc;
aud[41316]=16'hd7eb;
aud[41317]=16'hd7db;
aud[41318]=16'hd7ca;
aud[41319]=16'hd7b9;
aud[41320]=16'hd7a9;
aud[41321]=16'hd798;
aud[41322]=16'hd787;
aud[41323]=16'hd777;
aud[41324]=16'hd766;
aud[41325]=16'hd756;
aud[41326]=16'hd745;
aud[41327]=16'hd734;
aud[41328]=16'hd724;
aud[41329]=16'hd713;
aud[41330]=16'hd703;
aud[41331]=16'hd6f2;
aud[41332]=16'hd6e2;
aud[41333]=16'hd6d2;
aud[41334]=16'hd6c1;
aud[41335]=16'hd6b1;
aud[41336]=16'hd6a0;
aud[41337]=16'hd690;
aud[41338]=16'hd680;
aud[41339]=16'hd66f;
aud[41340]=16'hd65f;
aud[41341]=16'hd64f;
aud[41342]=16'hd63f;
aud[41343]=16'hd62e;
aud[41344]=16'hd61e;
aud[41345]=16'hd60e;
aud[41346]=16'hd5fe;
aud[41347]=16'hd5ee;
aud[41348]=16'hd5dd;
aud[41349]=16'hd5cd;
aud[41350]=16'hd5bd;
aud[41351]=16'hd5ad;
aud[41352]=16'hd59d;
aud[41353]=16'hd58d;
aud[41354]=16'hd57d;
aud[41355]=16'hd56d;
aud[41356]=16'hd55d;
aud[41357]=16'hd54d;
aud[41358]=16'hd53d;
aud[41359]=16'hd52d;
aud[41360]=16'hd51d;
aud[41361]=16'hd50d;
aud[41362]=16'hd4fd;
aud[41363]=16'hd4ed;
aud[41364]=16'hd4de;
aud[41365]=16'hd4ce;
aud[41366]=16'hd4be;
aud[41367]=16'hd4ae;
aud[41368]=16'hd49e;
aud[41369]=16'hd48f;
aud[41370]=16'hd47f;
aud[41371]=16'hd46f;
aud[41372]=16'hd45f;
aud[41373]=16'hd450;
aud[41374]=16'hd440;
aud[41375]=16'hd430;
aud[41376]=16'hd421;
aud[41377]=16'hd411;
aud[41378]=16'hd402;
aud[41379]=16'hd3f2;
aud[41380]=16'hd3e2;
aud[41381]=16'hd3d3;
aud[41382]=16'hd3c3;
aud[41383]=16'hd3b4;
aud[41384]=16'hd3a4;
aud[41385]=16'hd395;
aud[41386]=16'hd386;
aud[41387]=16'hd376;
aud[41388]=16'hd367;
aud[41389]=16'hd357;
aud[41390]=16'hd348;
aud[41391]=16'hd339;
aud[41392]=16'hd329;
aud[41393]=16'hd31a;
aud[41394]=16'hd30b;
aud[41395]=16'hd2fc;
aud[41396]=16'hd2ec;
aud[41397]=16'hd2dd;
aud[41398]=16'hd2ce;
aud[41399]=16'hd2bf;
aud[41400]=16'hd2b0;
aud[41401]=16'hd2a0;
aud[41402]=16'hd291;
aud[41403]=16'hd282;
aud[41404]=16'hd273;
aud[41405]=16'hd264;
aud[41406]=16'hd255;
aud[41407]=16'hd246;
aud[41408]=16'hd237;
aud[41409]=16'hd228;
aud[41410]=16'hd219;
aud[41411]=16'hd20a;
aud[41412]=16'hd1fb;
aud[41413]=16'hd1ec;
aud[41414]=16'hd1de;
aud[41415]=16'hd1cf;
aud[41416]=16'hd1c0;
aud[41417]=16'hd1b1;
aud[41418]=16'hd1a2;
aud[41419]=16'hd193;
aud[41420]=16'hd185;
aud[41421]=16'hd176;
aud[41422]=16'hd167;
aud[41423]=16'hd159;
aud[41424]=16'hd14a;
aud[41425]=16'hd13b;
aud[41426]=16'hd12d;
aud[41427]=16'hd11e;
aud[41428]=16'hd10f;
aud[41429]=16'hd101;
aud[41430]=16'hd0f2;
aud[41431]=16'hd0e4;
aud[41432]=16'hd0d5;
aud[41433]=16'hd0c7;
aud[41434]=16'hd0b8;
aud[41435]=16'hd0aa;
aud[41436]=16'hd09b;
aud[41437]=16'hd08d;
aud[41438]=16'hd07f;
aud[41439]=16'hd070;
aud[41440]=16'hd062;
aud[41441]=16'hd054;
aud[41442]=16'hd045;
aud[41443]=16'hd037;
aud[41444]=16'hd029;
aud[41445]=16'hd01b;
aud[41446]=16'hd00c;
aud[41447]=16'hcffe;
aud[41448]=16'hcff0;
aud[41449]=16'hcfe2;
aud[41450]=16'hcfd4;
aud[41451]=16'hcfc6;
aud[41452]=16'hcfb8;
aud[41453]=16'hcfa9;
aud[41454]=16'hcf9b;
aud[41455]=16'hcf8d;
aud[41456]=16'hcf7f;
aud[41457]=16'hcf71;
aud[41458]=16'hcf63;
aud[41459]=16'hcf56;
aud[41460]=16'hcf48;
aud[41461]=16'hcf3a;
aud[41462]=16'hcf2c;
aud[41463]=16'hcf1e;
aud[41464]=16'hcf10;
aud[41465]=16'hcf02;
aud[41466]=16'hcef5;
aud[41467]=16'hcee7;
aud[41468]=16'hced9;
aud[41469]=16'hcecb;
aud[41470]=16'hcebe;
aud[41471]=16'hceb0;
aud[41472]=16'hcea2;
aud[41473]=16'hce95;
aud[41474]=16'hce87;
aud[41475]=16'hce79;
aud[41476]=16'hce6c;
aud[41477]=16'hce5e;
aud[41478]=16'hce51;
aud[41479]=16'hce43;
aud[41480]=16'hce36;
aud[41481]=16'hce28;
aud[41482]=16'hce1b;
aud[41483]=16'hce0d;
aud[41484]=16'hce00;
aud[41485]=16'hcdf3;
aud[41486]=16'hcde5;
aud[41487]=16'hcdd8;
aud[41488]=16'hcdcb;
aud[41489]=16'hcdbd;
aud[41490]=16'hcdb0;
aud[41491]=16'hcda3;
aud[41492]=16'hcd96;
aud[41493]=16'hcd88;
aud[41494]=16'hcd7b;
aud[41495]=16'hcd6e;
aud[41496]=16'hcd61;
aud[41497]=16'hcd54;
aud[41498]=16'hcd47;
aud[41499]=16'hcd3a;
aud[41500]=16'hcd2d;
aud[41501]=16'hcd20;
aud[41502]=16'hcd13;
aud[41503]=16'hcd06;
aud[41504]=16'hccf9;
aud[41505]=16'hccec;
aud[41506]=16'hccdf;
aud[41507]=16'hccd2;
aud[41508]=16'hccc5;
aud[41509]=16'hccb8;
aud[41510]=16'hccab;
aud[41511]=16'hcc9f;
aud[41512]=16'hcc92;
aud[41513]=16'hcc85;
aud[41514]=16'hcc78;
aud[41515]=16'hcc6c;
aud[41516]=16'hcc5f;
aud[41517]=16'hcc52;
aud[41518]=16'hcc46;
aud[41519]=16'hcc39;
aud[41520]=16'hcc2c;
aud[41521]=16'hcc20;
aud[41522]=16'hcc13;
aud[41523]=16'hcc07;
aud[41524]=16'hcbfa;
aud[41525]=16'hcbee;
aud[41526]=16'hcbe1;
aud[41527]=16'hcbd5;
aud[41528]=16'hcbc9;
aud[41529]=16'hcbbc;
aud[41530]=16'hcbb0;
aud[41531]=16'hcba3;
aud[41532]=16'hcb97;
aud[41533]=16'hcb8b;
aud[41534]=16'hcb7f;
aud[41535]=16'hcb72;
aud[41536]=16'hcb66;
aud[41537]=16'hcb5a;
aud[41538]=16'hcb4e;
aud[41539]=16'hcb42;
aud[41540]=16'hcb35;
aud[41541]=16'hcb29;
aud[41542]=16'hcb1d;
aud[41543]=16'hcb11;
aud[41544]=16'hcb05;
aud[41545]=16'hcaf9;
aud[41546]=16'hcaed;
aud[41547]=16'hcae1;
aud[41548]=16'hcad5;
aud[41549]=16'hcac9;
aud[41550]=16'hcabd;
aud[41551]=16'hcab1;
aud[41552]=16'hcaa6;
aud[41553]=16'hca9a;
aud[41554]=16'hca8e;
aud[41555]=16'hca82;
aud[41556]=16'hca76;
aud[41557]=16'hca6b;
aud[41558]=16'hca5f;
aud[41559]=16'hca53;
aud[41560]=16'hca48;
aud[41561]=16'hca3c;
aud[41562]=16'hca30;
aud[41563]=16'hca25;
aud[41564]=16'hca19;
aud[41565]=16'hca0e;
aud[41566]=16'hca02;
aud[41567]=16'hc9f7;
aud[41568]=16'hc9eb;
aud[41569]=16'hc9e0;
aud[41570]=16'hc9d4;
aud[41571]=16'hc9c9;
aud[41572]=16'hc9bd;
aud[41573]=16'hc9b2;
aud[41574]=16'hc9a7;
aud[41575]=16'hc99b;
aud[41576]=16'hc990;
aud[41577]=16'hc985;
aud[41578]=16'hc97a;
aud[41579]=16'hc96e;
aud[41580]=16'hc963;
aud[41581]=16'hc958;
aud[41582]=16'hc94d;
aud[41583]=16'hc942;
aud[41584]=16'hc937;
aud[41585]=16'hc92c;
aud[41586]=16'hc920;
aud[41587]=16'hc915;
aud[41588]=16'hc90a;
aud[41589]=16'hc8ff;
aud[41590]=16'hc8f5;
aud[41591]=16'hc8ea;
aud[41592]=16'hc8df;
aud[41593]=16'hc8d4;
aud[41594]=16'hc8c9;
aud[41595]=16'hc8be;
aud[41596]=16'hc8b3;
aud[41597]=16'hc8a9;
aud[41598]=16'hc89e;
aud[41599]=16'hc893;
aud[41600]=16'hc888;
aud[41601]=16'hc87e;
aud[41602]=16'hc873;
aud[41603]=16'hc868;
aud[41604]=16'hc85e;
aud[41605]=16'hc853;
aud[41606]=16'hc849;
aud[41607]=16'hc83e;
aud[41608]=16'hc834;
aud[41609]=16'hc829;
aud[41610]=16'hc81f;
aud[41611]=16'hc814;
aud[41612]=16'hc80a;
aud[41613]=16'hc7ff;
aud[41614]=16'hc7f5;
aud[41615]=16'hc7eb;
aud[41616]=16'hc7e0;
aud[41617]=16'hc7d6;
aud[41618]=16'hc7cc;
aud[41619]=16'hc7c1;
aud[41620]=16'hc7b7;
aud[41621]=16'hc7ad;
aud[41622]=16'hc7a3;
aud[41623]=16'hc799;
aud[41624]=16'hc78f;
aud[41625]=16'hc785;
aud[41626]=16'hc77a;
aud[41627]=16'hc770;
aud[41628]=16'hc766;
aud[41629]=16'hc75c;
aud[41630]=16'hc752;
aud[41631]=16'hc748;
aud[41632]=16'hc73f;
aud[41633]=16'hc735;
aud[41634]=16'hc72b;
aud[41635]=16'hc721;
aud[41636]=16'hc717;
aud[41637]=16'hc70d;
aud[41638]=16'hc703;
aud[41639]=16'hc6fa;
aud[41640]=16'hc6f0;
aud[41641]=16'hc6e6;
aud[41642]=16'hc6dd;
aud[41643]=16'hc6d3;
aud[41644]=16'hc6c9;
aud[41645]=16'hc6c0;
aud[41646]=16'hc6b6;
aud[41647]=16'hc6ad;
aud[41648]=16'hc6a3;
aud[41649]=16'hc69a;
aud[41650]=16'hc690;
aud[41651]=16'hc687;
aud[41652]=16'hc67d;
aud[41653]=16'hc674;
aud[41654]=16'hc66b;
aud[41655]=16'hc661;
aud[41656]=16'hc658;
aud[41657]=16'hc64f;
aud[41658]=16'hc645;
aud[41659]=16'hc63c;
aud[41660]=16'hc633;
aud[41661]=16'hc62a;
aud[41662]=16'hc620;
aud[41663]=16'hc617;
aud[41664]=16'hc60e;
aud[41665]=16'hc605;
aud[41666]=16'hc5fc;
aud[41667]=16'hc5f3;
aud[41668]=16'hc5ea;
aud[41669]=16'hc5e1;
aud[41670]=16'hc5d8;
aud[41671]=16'hc5cf;
aud[41672]=16'hc5c6;
aud[41673]=16'hc5bd;
aud[41674]=16'hc5b4;
aud[41675]=16'hc5ac;
aud[41676]=16'hc5a3;
aud[41677]=16'hc59a;
aud[41678]=16'hc591;
aud[41679]=16'hc588;
aud[41680]=16'hc580;
aud[41681]=16'hc577;
aud[41682]=16'hc56e;
aud[41683]=16'hc566;
aud[41684]=16'hc55d;
aud[41685]=16'hc555;
aud[41686]=16'hc54c;
aud[41687]=16'hc544;
aud[41688]=16'hc53b;
aud[41689]=16'hc533;
aud[41690]=16'hc52a;
aud[41691]=16'hc522;
aud[41692]=16'hc519;
aud[41693]=16'hc511;
aud[41694]=16'hc509;
aud[41695]=16'hc500;
aud[41696]=16'hc4f8;
aud[41697]=16'hc4f0;
aud[41698]=16'hc4e7;
aud[41699]=16'hc4df;
aud[41700]=16'hc4d7;
aud[41701]=16'hc4cf;
aud[41702]=16'hc4c7;
aud[41703]=16'hc4bf;
aud[41704]=16'hc4b6;
aud[41705]=16'hc4ae;
aud[41706]=16'hc4a6;
aud[41707]=16'hc49e;
aud[41708]=16'hc496;
aud[41709]=16'hc48e;
aud[41710]=16'hc486;
aud[41711]=16'hc47f;
aud[41712]=16'hc477;
aud[41713]=16'hc46f;
aud[41714]=16'hc467;
aud[41715]=16'hc45f;
aud[41716]=16'hc457;
aud[41717]=16'hc450;
aud[41718]=16'hc448;
aud[41719]=16'hc440;
aud[41720]=16'hc439;
aud[41721]=16'hc431;
aud[41722]=16'hc429;
aud[41723]=16'hc422;
aud[41724]=16'hc41a;
aud[41725]=16'hc413;
aud[41726]=16'hc40b;
aud[41727]=16'hc404;
aud[41728]=16'hc3fc;
aud[41729]=16'hc3f5;
aud[41730]=16'hc3ed;
aud[41731]=16'hc3e6;
aud[41732]=16'hc3df;
aud[41733]=16'hc3d7;
aud[41734]=16'hc3d0;
aud[41735]=16'hc3c9;
aud[41736]=16'hc3c1;
aud[41737]=16'hc3ba;
aud[41738]=16'hc3b3;
aud[41739]=16'hc3ac;
aud[41740]=16'hc3a5;
aud[41741]=16'hc39d;
aud[41742]=16'hc396;
aud[41743]=16'hc38f;
aud[41744]=16'hc388;
aud[41745]=16'hc381;
aud[41746]=16'hc37a;
aud[41747]=16'hc373;
aud[41748]=16'hc36c;
aud[41749]=16'hc365;
aud[41750]=16'hc35f;
aud[41751]=16'hc358;
aud[41752]=16'hc351;
aud[41753]=16'hc34a;
aud[41754]=16'hc343;
aud[41755]=16'hc33d;
aud[41756]=16'hc336;
aud[41757]=16'hc32f;
aud[41758]=16'hc329;
aud[41759]=16'hc322;
aud[41760]=16'hc31b;
aud[41761]=16'hc315;
aud[41762]=16'hc30e;
aud[41763]=16'hc308;
aud[41764]=16'hc301;
aud[41765]=16'hc2fb;
aud[41766]=16'hc2f4;
aud[41767]=16'hc2ee;
aud[41768]=16'hc2e7;
aud[41769]=16'hc2e1;
aud[41770]=16'hc2db;
aud[41771]=16'hc2d4;
aud[41772]=16'hc2ce;
aud[41773]=16'hc2c8;
aud[41774]=16'hc2c1;
aud[41775]=16'hc2bb;
aud[41776]=16'hc2b5;
aud[41777]=16'hc2af;
aud[41778]=16'hc2a9;
aud[41779]=16'hc2a3;
aud[41780]=16'hc29d;
aud[41781]=16'hc297;
aud[41782]=16'hc291;
aud[41783]=16'hc28b;
aud[41784]=16'hc285;
aud[41785]=16'hc27f;
aud[41786]=16'hc279;
aud[41787]=16'hc273;
aud[41788]=16'hc26d;
aud[41789]=16'hc267;
aud[41790]=16'hc261;
aud[41791]=16'hc25c;
aud[41792]=16'hc256;
aud[41793]=16'hc250;
aud[41794]=16'hc24a;
aud[41795]=16'hc245;
aud[41796]=16'hc23f;
aud[41797]=16'hc239;
aud[41798]=16'hc234;
aud[41799]=16'hc22e;
aud[41800]=16'hc229;
aud[41801]=16'hc223;
aud[41802]=16'hc21e;
aud[41803]=16'hc218;
aud[41804]=16'hc213;
aud[41805]=16'hc20d;
aud[41806]=16'hc208;
aud[41807]=16'hc203;
aud[41808]=16'hc1fd;
aud[41809]=16'hc1f8;
aud[41810]=16'hc1f3;
aud[41811]=16'hc1ee;
aud[41812]=16'hc1e8;
aud[41813]=16'hc1e3;
aud[41814]=16'hc1de;
aud[41815]=16'hc1d9;
aud[41816]=16'hc1d4;
aud[41817]=16'hc1cf;
aud[41818]=16'hc1ca;
aud[41819]=16'hc1c5;
aud[41820]=16'hc1c0;
aud[41821]=16'hc1bb;
aud[41822]=16'hc1b6;
aud[41823]=16'hc1b1;
aud[41824]=16'hc1ac;
aud[41825]=16'hc1a7;
aud[41826]=16'hc1a2;
aud[41827]=16'hc19e;
aud[41828]=16'hc199;
aud[41829]=16'hc194;
aud[41830]=16'hc18f;
aud[41831]=16'hc18b;
aud[41832]=16'hc186;
aud[41833]=16'hc181;
aud[41834]=16'hc17d;
aud[41835]=16'hc178;
aud[41836]=16'hc174;
aud[41837]=16'hc16f;
aud[41838]=16'hc16b;
aud[41839]=16'hc166;
aud[41840]=16'hc162;
aud[41841]=16'hc15d;
aud[41842]=16'hc159;
aud[41843]=16'hc154;
aud[41844]=16'hc150;
aud[41845]=16'hc14c;
aud[41846]=16'hc147;
aud[41847]=16'hc143;
aud[41848]=16'hc13f;
aud[41849]=16'hc13b;
aud[41850]=16'hc137;
aud[41851]=16'hc133;
aud[41852]=16'hc12e;
aud[41853]=16'hc12a;
aud[41854]=16'hc126;
aud[41855]=16'hc122;
aud[41856]=16'hc11e;
aud[41857]=16'hc11a;
aud[41858]=16'hc116;
aud[41859]=16'hc112;
aud[41860]=16'hc10e;
aud[41861]=16'hc10b;
aud[41862]=16'hc107;
aud[41863]=16'hc103;
aud[41864]=16'hc0ff;
aud[41865]=16'hc0fb;
aud[41866]=16'hc0f8;
aud[41867]=16'hc0f4;
aud[41868]=16'hc0f0;
aud[41869]=16'hc0ed;
aud[41870]=16'hc0e9;
aud[41871]=16'hc0e5;
aud[41872]=16'hc0e2;
aud[41873]=16'hc0de;
aud[41874]=16'hc0db;
aud[41875]=16'hc0d7;
aud[41876]=16'hc0d4;
aud[41877]=16'hc0d0;
aud[41878]=16'hc0cd;
aud[41879]=16'hc0ca;
aud[41880]=16'hc0c6;
aud[41881]=16'hc0c3;
aud[41882]=16'hc0c0;
aud[41883]=16'hc0bd;
aud[41884]=16'hc0b9;
aud[41885]=16'hc0b6;
aud[41886]=16'hc0b3;
aud[41887]=16'hc0b0;
aud[41888]=16'hc0ad;
aud[41889]=16'hc0aa;
aud[41890]=16'hc0a6;
aud[41891]=16'hc0a3;
aud[41892]=16'hc0a0;
aud[41893]=16'hc09d;
aud[41894]=16'hc09b;
aud[41895]=16'hc098;
aud[41896]=16'hc095;
aud[41897]=16'hc092;
aud[41898]=16'hc08f;
aud[41899]=16'hc08c;
aud[41900]=16'hc089;
aud[41901]=16'hc087;
aud[41902]=16'hc084;
aud[41903]=16'hc081;
aud[41904]=16'hc07f;
aud[41905]=16'hc07c;
aud[41906]=16'hc079;
aud[41907]=16'hc077;
aud[41908]=16'hc074;
aud[41909]=16'hc072;
aud[41910]=16'hc06f;
aud[41911]=16'hc06d;
aud[41912]=16'hc06a;
aud[41913]=16'hc068;
aud[41914]=16'hc065;
aud[41915]=16'hc063;
aud[41916]=16'hc061;
aud[41917]=16'hc05e;
aud[41918]=16'hc05c;
aud[41919]=16'hc05a;
aud[41920]=16'hc058;
aud[41921]=16'hc055;
aud[41922]=16'hc053;
aud[41923]=16'hc051;
aud[41924]=16'hc04f;
aud[41925]=16'hc04d;
aud[41926]=16'hc04b;
aud[41927]=16'hc049;
aud[41928]=16'hc047;
aud[41929]=16'hc045;
aud[41930]=16'hc043;
aud[41931]=16'hc041;
aud[41932]=16'hc03f;
aud[41933]=16'hc03d;
aud[41934]=16'hc03b;
aud[41935]=16'hc039;
aud[41936]=16'hc038;
aud[41937]=16'hc036;
aud[41938]=16'hc034;
aud[41939]=16'hc033;
aud[41940]=16'hc031;
aud[41941]=16'hc02f;
aud[41942]=16'hc02e;
aud[41943]=16'hc02c;
aud[41944]=16'hc02a;
aud[41945]=16'hc029;
aud[41946]=16'hc027;
aud[41947]=16'hc026;
aud[41948]=16'hc024;
aud[41949]=16'hc023;
aud[41950]=16'hc022;
aud[41951]=16'hc020;
aud[41952]=16'hc01f;
aud[41953]=16'hc01e;
aud[41954]=16'hc01c;
aud[41955]=16'hc01b;
aud[41956]=16'hc01a;
aud[41957]=16'hc019;
aud[41958]=16'hc018;
aud[41959]=16'hc016;
aud[41960]=16'hc015;
aud[41961]=16'hc014;
aud[41962]=16'hc013;
aud[41963]=16'hc012;
aud[41964]=16'hc011;
aud[41965]=16'hc010;
aud[41966]=16'hc00f;
aud[41967]=16'hc00e;
aud[41968]=16'hc00d;
aud[41969]=16'hc00d;
aud[41970]=16'hc00c;
aud[41971]=16'hc00b;
aud[41972]=16'hc00a;
aud[41973]=16'hc009;
aud[41974]=16'hc009;
aud[41975]=16'hc008;
aud[41976]=16'hc007;
aud[41977]=16'hc007;
aud[41978]=16'hc006;
aud[41979]=16'hc006;
aud[41980]=16'hc005;
aud[41981]=16'hc005;
aud[41982]=16'hc004;
aud[41983]=16'hc004;
aud[41984]=16'hc003;
aud[41985]=16'hc003;
aud[41986]=16'hc002;
aud[41987]=16'hc002;
aud[41988]=16'hc002;
aud[41989]=16'hc001;
aud[41990]=16'hc001;
aud[41991]=16'hc001;
aud[41992]=16'hc001;
aud[41993]=16'hc001;
aud[41994]=16'hc000;
aud[41995]=16'hc000;
aud[41996]=16'hc000;
aud[41997]=16'hc000;
aud[41998]=16'hc000;
aud[41999]=16'hc000;
aud[42000]=16'hc000;
aud[42001]=16'hc000;
aud[42002]=16'hc000;
aud[42003]=16'hc000;
aud[42004]=16'hc000;
aud[42005]=16'hc001;
aud[42006]=16'hc001;
aud[42007]=16'hc001;
aud[42008]=16'hc001;
aud[42009]=16'hc001;
aud[42010]=16'hc002;
aud[42011]=16'hc002;
aud[42012]=16'hc002;
aud[42013]=16'hc003;
aud[42014]=16'hc003;
aud[42015]=16'hc004;
aud[42016]=16'hc004;
aud[42017]=16'hc005;
aud[42018]=16'hc005;
aud[42019]=16'hc006;
aud[42020]=16'hc006;
aud[42021]=16'hc007;
aud[42022]=16'hc007;
aud[42023]=16'hc008;
aud[42024]=16'hc009;
aud[42025]=16'hc009;
aud[42026]=16'hc00a;
aud[42027]=16'hc00b;
aud[42028]=16'hc00c;
aud[42029]=16'hc00d;
aud[42030]=16'hc00d;
aud[42031]=16'hc00e;
aud[42032]=16'hc00f;
aud[42033]=16'hc010;
aud[42034]=16'hc011;
aud[42035]=16'hc012;
aud[42036]=16'hc013;
aud[42037]=16'hc014;
aud[42038]=16'hc015;
aud[42039]=16'hc016;
aud[42040]=16'hc018;
aud[42041]=16'hc019;
aud[42042]=16'hc01a;
aud[42043]=16'hc01b;
aud[42044]=16'hc01c;
aud[42045]=16'hc01e;
aud[42046]=16'hc01f;
aud[42047]=16'hc020;
aud[42048]=16'hc022;
aud[42049]=16'hc023;
aud[42050]=16'hc024;
aud[42051]=16'hc026;
aud[42052]=16'hc027;
aud[42053]=16'hc029;
aud[42054]=16'hc02a;
aud[42055]=16'hc02c;
aud[42056]=16'hc02e;
aud[42057]=16'hc02f;
aud[42058]=16'hc031;
aud[42059]=16'hc033;
aud[42060]=16'hc034;
aud[42061]=16'hc036;
aud[42062]=16'hc038;
aud[42063]=16'hc039;
aud[42064]=16'hc03b;
aud[42065]=16'hc03d;
aud[42066]=16'hc03f;
aud[42067]=16'hc041;
aud[42068]=16'hc043;
aud[42069]=16'hc045;
aud[42070]=16'hc047;
aud[42071]=16'hc049;
aud[42072]=16'hc04b;
aud[42073]=16'hc04d;
aud[42074]=16'hc04f;
aud[42075]=16'hc051;
aud[42076]=16'hc053;
aud[42077]=16'hc055;
aud[42078]=16'hc058;
aud[42079]=16'hc05a;
aud[42080]=16'hc05c;
aud[42081]=16'hc05e;
aud[42082]=16'hc061;
aud[42083]=16'hc063;
aud[42084]=16'hc065;
aud[42085]=16'hc068;
aud[42086]=16'hc06a;
aud[42087]=16'hc06d;
aud[42088]=16'hc06f;
aud[42089]=16'hc072;
aud[42090]=16'hc074;
aud[42091]=16'hc077;
aud[42092]=16'hc079;
aud[42093]=16'hc07c;
aud[42094]=16'hc07f;
aud[42095]=16'hc081;
aud[42096]=16'hc084;
aud[42097]=16'hc087;
aud[42098]=16'hc089;
aud[42099]=16'hc08c;
aud[42100]=16'hc08f;
aud[42101]=16'hc092;
aud[42102]=16'hc095;
aud[42103]=16'hc098;
aud[42104]=16'hc09b;
aud[42105]=16'hc09d;
aud[42106]=16'hc0a0;
aud[42107]=16'hc0a3;
aud[42108]=16'hc0a6;
aud[42109]=16'hc0aa;
aud[42110]=16'hc0ad;
aud[42111]=16'hc0b0;
aud[42112]=16'hc0b3;
aud[42113]=16'hc0b6;
aud[42114]=16'hc0b9;
aud[42115]=16'hc0bd;
aud[42116]=16'hc0c0;
aud[42117]=16'hc0c3;
aud[42118]=16'hc0c6;
aud[42119]=16'hc0ca;
aud[42120]=16'hc0cd;
aud[42121]=16'hc0d0;
aud[42122]=16'hc0d4;
aud[42123]=16'hc0d7;
aud[42124]=16'hc0db;
aud[42125]=16'hc0de;
aud[42126]=16'hc0e2;
aud[42127]=16'hc0e5;
aud[42128]=16'hc0e9;
aud[42129]=16'hc0ed;
aud[42130]=16'hc0f0;
aud[42131]=16'hc0f4;
aud[42132]=16'hc0f8;
aud[42133]=16'hc0fb;
aud[42134]=16'hc0ff;
aud[42135]=16'hc103;
aud[42136]=16'hc107;
aud[42137]=16'hc10b;
aud[42138]=16'hc10e;
aud[42139]=16'hc112;
aud[42140]=16'hc116;
aud[42141]=16'hc11a;
aud[42142]=16'hc11e;
aud[42143]=16'hc122;
aud[42144]=16'hc126;
aud[42145]=16'hc12a;
aud[42146]=16'hc12e;
aud[42147]=16'hc133;
aud[42148]=16'hc137;
aud[42149]=16'hc13b;
aud[42150]=16'hc13f;
aud[42151]=16'hc143;
aud[42152]=16'hc147;
aud[42153]=16'hc14c;
aud[42154]=16'hc150;
aud[42155]=16'hc154;
aud[42156]=16'hc159;
aud[42157]=16'hc15d;
aud[42158]=16'hc162;
aud[42159]=16'hc166;
aud[42160]=16'hc16b;
aud[42161]=16'hc16f;
aud[42162]=16'hc174;
aud[42163]=16'hc178;
aud[42164]=16'hc17d;
aud[42165]=16'hc181;
aud[42166]=16'hc186;
aud[42167]=16'hc18b;
aud[42168]=16'hc18f;
aud[42169]=16'hc194;
aud[42170]=16'hc199;
aud[42171]=16'hc19e;
aud[42172]=16'hc1a2;
aud[42173]=16'hc1a7;
aud[42174]=16'hc1ac;
aud[42175]=16'hc1b1;
aud[42176]=16'hc1b6;
aud[42177]=16'hc1bb;
aud[42178]=16'hc1c0;
aud[42179]=16'hc1c5;
aud[42180]=16'hc1ca;
aud[42181]=16'hc1cf;
aud[42182]=16'hc1d4;
aud[42183]=16'hc1d9;
aud[42184]=16'hc1de;
aud[42185]=16'hc1e3;
aud[42186]=16'hc1e8;
aud[42187]=16'hc1ee;
aud[42188]=16'hc1f3;
aud[42189]=16'hc1f8;
aud[42190]=16'hc1fd;
aud[42191]=16'hc203;
aud[42192]=16'hc208;
aud[42193]=16'hc20d;
aud[42194]=16'hc213;
aud[42195]=16'hc218;
aud[42196]=16'hc21e;
aud[42197]=16'hc223;
aud[42198]=16'hc229;
aud[42199]=16'hc22e;
aud[42200]=16'hc234;
aud[42201]=16'hc239;
aud[42202]=16'hc23f;
aud[42203]=16'hc245;
aud[42204]=16'hc24a;
aud[42205]=16'hc250;
aud[42206]=16'hc256;
aud[42207]=16'hc25c;
aud[42208]=16'hc261;
aud[42209]=16'hc267;
aud[42210]=16'hc26d;
aud[42211]=16'hc273;
aud[42212]=16'hc279;
aud[42213]=16'hc27f;
aud[42214]=16'hc285;
aud[42215]=16'hc28b;
aud[42216]=16'hc291;
aud[42217]=16'hc297;
aud[42218]=16'hc29d;
aud[42219]=16'hc2a3;
aud[42220]=16'hc2a9;
aud[42221]=16'hc2af;
aud[42222]=16'hc2b5;
aud[42223]=16'hc2bb;
aud[42224]=16'hc2c1;
aud[42225]=16'hc2c8;
aud[42226]=16'hc2ce;
aud[42227]=16'hc2d4;
aud[42228]=16'hc2db;
aud[42229]=16'hc2e1;
aud[42230]=16'hc2e7;
aud[42231]=16'hc2ee;
aud[42232]=16'hc2f4;
aud[42233]=16'hc2fb;
aud[42234]=16'hc301;
aud[42235]=16'hc308;
aud[42236]=16'hc30e;
aud[42237]=16'hc315;
aud[42238]=16'hc31b;
aud[42239]=16'hc322;
aud[42240]=16'hc329;
aud[42241]=16'hc32f;
aud[42242]=16'hc336;
aud[42243]=16'hc33d;
aud[42244]=16'hc343;
aud[42245]=16'hc34a;
aud[42246]=16'hc351;
aud[42247]=16'hc358;
aud[42248]=16'hc35f;
aud[42249]=16'hc365;
aud[42250]=16'hc36c;
aud[42251]=16'hc373;
aud[42252]=16'hc37a;
aud[42253]=16'hc381;
aud[42254]=16'hc388;
aud[42255]=16'hc38f;
aud[42256]=16'hc396;
aud[42257]=16'hc39d;
aud[42258]=16'hc3a5;
aud[42259]=16'hc3ac;
aud[42260]=16'hc3b3;
aud[42261]=16'hc3ba;
aud[42262]=16'hc3c1;
aud[42263]=16'hc3c9;
aud[42264]=16'hc3d0;
aud[42265]=16'hc3d7;
aud[42266]=16'hc3df;
aud[42267]=16'hc3e6;
aud[42268]=16'hc3ed;
aud[42269]=16'hc3f5;
aud[42270]=16'hc3fc;
aud[42271]=16'hc404;
aud[42272]=16'hc40b;
aud[42273]=16'hc413;
aud[42274]=16'hc41a;
aud[42275]=16'hc422;
aud[42276]=16'hc429;
aud[42277]=16'hc431;
aud[42278]=16'hc439;
aud[42279]=16'hc440;
aud[42280]=16'hc448;
aud[42281]=16'hc450;
aud[42282]=16'hc457;
aud[42283]=16'hc45f;
aud[42284]=16'hc467;
aud[42285]=16'hc46f;
aud[42286]=16'hc477;
aud[42287]=16'hc47f;
aud[42288]=16'hc486;
aud[42289]=16'hc48e;
aud[42290]=16'hc496;
aud[42291]=16'hc49e;
aud[42292]=16'hc4a6;
aud[42293]=16'hc4ae;
aud[42294]=16'hc4b6;
aud[42295]=16'hc4bf;
aud[42296]=16'hc4c7;
aud[42297]=16'hc4cf;
aud[42298]=16'hc4d7;
aud[42299]=16'hc4df;
aud[42300]=16'hc4e7;
aud[42301]=16'hc4f0;
aud[42302]=16'hc4f8;
aud[42303]=16'hc500;
aud[42304]=16'hc509;
aud[42305]=16'hc511;
aud[42306]=16'hc519;
aud[42307]=16'hc522;
aud[42308]=16'hc52a;
aud[42309]=16'hc533;
aud[42310]=16'hc53b;
aud[42311]=16'hc544;
aud[42312]=16'hc54c;
aud[42313]=16'hc555;
aud[42314]=16'hc55d;
aud[42315]=16'hc566;
aud[42316]=16'hc56e;
aud[42317]=16'hc577;
aud[42318]=16'hc580;
aud[42319]=16'hc588;
aud[42320]=16'hc591;
aud[42321]=16'hc59a;
aud[42322]=16'hc5a3;
aud[42323]=16'hc5ac;
aud[42324]=16'hc5b4;
aud[42325]=16'hc5bd;
aud[42326]=16'hc5c6;
aud[42327]=16'hc5cf;
aud[42328]=16'hc5d8;
aud[42329]=16'hc5e1;
aud[42330]=16'hc5ea;
aud[42331]=16'hc5f3;
aud[42332]=16'hc5fc;
aud[42333]=16'hc605;
aud[42334]=16'hc60e;
aud[42335]=16'hc617;
aud[42336]=16'hc620;
aud[42337]=16'hc62a;
aud[42338]=16'hc633;
aud[42339]=16'hc63c;
aud[42340]=16'hc645;
aud[42341]=16'hc64f;
aud[42342]=16'hc658;
aud[42343]=16'hc661;
aud[42344]=16'hc66b;
aud[42345]=16'hc674;
aud[42346]=16'hc67d;
aud[42347]=16'hc687;
aud[42348]=16'hc690;
aud[42349]=16'hc69a;
aud[42350]=16'hc6a3;
aud[42351]=16'hc6ad;
aud[42352]=16'hc6b6;
aud[42353]=16'hc6c0;
aud[42354]=16'hc6c9;
aud[42355]=16'hc6d3;
aud[42356]=16'hc6dd;
aud[42357]=16'hc6e6;
aud[42358]=16'hc6f0;
aud[42359]=16'hc6fa;
aud[42360]=16'hc703;
aud[42361]=16'hc70d;
aud[42362]=16'hc717;
aud[42363]=16'hc721;
aud[42364]=16'hc72b;
aud[42365]=16'hc735;
aud[42366]=16'hc73f;
aud[42367]=16'hc748;
aud[42368]=16'hc752;
aud[42369]=16'hc75c;
aud[42370]=16'hc766;
aud[42371]=16'hc770;
aud[42372]=16'hc77a;
aud[42373]=16'hc785;
aud[42374]=16'hc78f;
aud[42375]=16'hc799;
aud[42376]=16'hc7a3;
aud[42377]=16'hc7ad;
aud[42378]=16'hc7b7;
aud[42379]=16'hc7c1;
aud[42380]=16'hc7cc;
aud[42381]=16'hc7d6;
aud[42382]=16'hc7e0;
aud[42383]=16'hc7eb;
aud[42384]=16'hc7f5;
aud[42385]=16'hc7ff;
aud[42386]=16'hc80a;
aud[42387]=16'hc814;
aud[42388]=16'hc81f;
aud[42389]=16'hc829;
aud[42390]=16'hc834;
aud[42391]=16'hc83e;
aud[42392]=16'hc849;
aud[42393]=16'hc853;
aud[42394]=16'hc85e;
aud[42395]=16'hc868;
aud[42396]=16'hc873;
aud[42397]=16'hc87e;
aud[42398]=16'hc888;
aud[42399]=16'hc893;
aud[42400]=16'hc89e;
aud[42401]=16'hc8a9;
aud[42402]=16'hc8b3;
aud[42403]=16'hc8be;
aud[42404]=16'hc8c9;
aud[42405]=16'hc8d4;
aud[42406]=16'hc8df;
aud[42407]=16'hc8ea;
aud[42408]=16'hc8f5;
aud[42409]=16'hc8ff;
aud[42410]=16'hc90a;
aud[42411]=16'hc915;
aud[42412]=16'hc920;
aud[42413]=16'hc92c;
aud[42414]=16'hc937;
aud[42415]=16'hc942;
aud[42416]=16'hc94d;
aud[42417]=16'hc958;
aud[42418]=16'hc963;
aud[42419]=16'hc96e;
aud[42420]=16'hc97a;
aud[42421]=16'hc985;
aud[42422]=16'hc990;
aud[42423]=16'hc99b;
aud[42424]=16'hc9a7;
aud[42425]=16'hc9b2;
aud[42426]=16'hc9bd;
aud[42427]=16'hc9c9;
aud[42428]=16'hc9d4;
aud[42429]=16'hc9e0;
aud[42430]=16'hc9eb;
aud[42431]=16'hc9f7;
aud[42432]=16'hca02;
aud[42433]=16'hca0e;
aud[42434]=16'hca19;
aud[42435]=16'hca25;
aud[42436]=16'hca30;
aud[42437]=16'hca3c;
aud[42438]=16'hca48;
aud[42439]=16'hca53;
aud[42440]=16'hca5f;
aud[42441]=16'hca6b;
aud[42442]=16'hca76;
aud[42443]=16'hca82;
aud[42444]=16'hca8e;
aud[42445]=16'hca9a;
aud[42446]=16'hcaa6;
aud[42447]=16'hcab1;
aud[42448]=16'hcabd;
aud[42449]=16'hcac9;
aud[42450]=16'hcad5;
aud[42451]=16'hcae1;
aud[42452]=16'hcaed;
aud[42453]=16'hcaf9;
aud[42454]=16'hcb05;
aud[42455]=16'hcb11;
aud[42456]=16'hcb1d;
aud[42457]=16'hcb29;
aud[42458]=16'hcb35;
aud[42459]=16'hcb42;
aud[42460]=16'hcb4e;
aud[42461]=16'hcb5a;
aud[42462]=16'hcb66;
aud[42463]=16'hcb72;
aud[42464]=16'hcb7f;
aud[42465]=16'hcb8b;
aud[42466]=16'hcb97;
aud[42467]=16'hcba3;
aud[42468]=16'hcbb0;
aud[42469]=16'hcbbc;
aud[42470]=16'hcbc9;
aud[42471]=16'hcbd5;
aud[42472]=16'hcbe1;
aud[42473]=16'hcbee;
aud[42474]=16'hcbfa;
aud[42475]=16'hcc07;
aud[42476]=16'hcc13;
aud[42477]=16'hcc20;
aud[42478]=16'hcc2c;
aud[42479]=16'hcc39;
aud[42480]=16'hcc46;
aud[42481]=16'hcc52;
aud[42482]=16'hcc5f;
aud[42483]=16'hcc6c;
aud[42484]=16'hcc78;
aud[42485]=16'hcc85;
aud[42486]=16'hcc92;
aud[42487]=16'hcc9f;
aud[42488]=16'hccab;
aud[42489]=16'hccb8;
aud[42490]=16'hccc5;
aud[42491]=16'hccd2;
aud[42492]=16'hccdf;
aud[42493]=16'hccec;
aud[42494]=16'hccf9;
aud[42495]=16'hcd06;
aud[42496]=16'hcd13;
aud[42497]=16'hcd20;
aud[42498]=16'hcd2d;
aud[42499]=16'hcd3a;
aud[42500]=16'hcd47;
aud[42501]=16'hcd54;
aud[42502]=16'hcd61;
aud[42503]=16'hcd6e;
aud[42504]=16'hcd7b;
aud[42505]=16'hcd88;
aud[42506]=16'hcd96;
aud[42507]=16'hcda3;
aud[42508]=16'hcdb0;
aud[42509]=16'hcdbd;
aud[42510]=16'hcdcb;
aud[42511]=16'hcdd8;
aud[42512]=16'hcde5;
aud[42513]=16'hcdf3;
aud[42514]=16'hce00;
aud[42515]=16'hce0d;
aud[42516]=16'hce1b;
aud[42517]=16'hce28;
aud[42518]=16'hce36;
aud[42519]=16'hce43;
aud[42520]=16'hce51;
aud[42521]=16'hce5e;
aud[42522]=16'hce6c;
aud[42523]=16'hce79;
aud[42524]=16'hce87;
aud[42525]=16'hce95;
aud[42526]=16'hcea2;
aud[42527]=16'hceb0;
aud[42528]=16'hcebe;
aud[42529]=16'hcecb;
aud[42530]=16'hced9;
aud[42531]=16'hcee7;
aud[42532]=16'hcef5;
aud[42533]=16'hcf02;
aud[42534]=16'hcf10;
aud[42535]=16'hcf1e;
aud[42536]=16'hcf2c;
aud[42537]=16'hcf3a;
aud[42538]=16'hcf48;
aud[42539]=16'hcf56;
aud[42540]=16'hcf63;
aud[42541]=16'hcf71;
aud[42542]=16'hcf7f;
aud[42543]=16'hcf8d;
aud[42544]=16'hcf9b;
aud[42545]=16'hcfa9;
aud[42546]=16'hcfb8;
aud[42547]=16'hcfc6;
aud[42548]=16'hcfd4;
aud[42549]=16'hcfe2;
aud[42550]=16'hcff0;
aud[42551]=16'hcffe;
aud[42552]=16'hd00c;
aud[42553]=16'hd01b;
aud[42554]=16'hd029;
aud[42555]=16'hd037;
aud[42556]=16'hd045;
aud[42557]=16'hd054;
aud[42558]=16'hd062;
aud[42559]=16'hd070;
aud[42560]=16'hd07f;
aud[42561]=16'hd08d;
aud[42562]=16'hd09b;
aud[42563]=16'hd0aa;
aud[42564]=16'hd0b8;
aud[42565]=16'hd0c7;
aud[42566]=16'hd0d5;
aud[42567]=16'hd0e4;
aud[42568]=16'hd0f2;
aud[42569]=16'hd101;
aud[42570]=16'hd10f;
aud[42571]=16'hd11e;
aud[42572]=16'hd12d;
aud[42573]=16'hd13b;
aud[42574]=16'hd14a;
aud[42575]=16'hd159;
aud[42576]=16'hd167;
aud[42577]=16'hd176;
aud[42578]=16'hd185;
aud[42579]=16'hd193;
aud[42580]=16'hd1a2;
aud[42581]=16'hd1b1;
aud[42582]=16'hd1c0;
aud[42583]=16'hd1cf;
aud[42584]=16'hd1de;
aud[42585]=16'hd1ec;
aud[42586]=16'hd1fb;
aud[42587]=16'hd20a;
aud[42588]=16'hd219;
aud[42589]=16'hd228;
aud[42590]=16'hd237;
aud[42591]=16'hd246;
aud[42592]=16'hd255;
aud[42593]=16'hd264;
aud[42594]=16'hd273;
aud[42595]=16'hd282;
aud[42596]=16'hd291;
aud[42597]=16'hd2a0;
aud[42598]=16'hd2b0;
aud[42599]=16'hd2bf;
aud[42600]=16'hd2ce;
aud[42601]=16'hd2dd;
aud[42602]=16'hd2ec;
aud[42603]=16'hd2fc;
aud[42604]=16'hd30b;
aud[42605]=16'hd31a;
aud[42606]=16'hd329;
aud[42607]=16'hd339;
aud[42608]=16'hd348;
aud[42609]=16'hd357;
aud[42610]=16'hd367;
aud[42611]=16'hd376;
aud[42612]=16'hd386;
aud[42613]=16'hd395;
aud[42614]=16'hd3a4;
aud[42615]=16'hd3b4;
aud[42616]=16'hd3c3;
aud[42617]=16'hd3d3;
aud[42618]=16'hd3e2;
aud[42619]=16'hd3f2;
aud[42620]=16'hd402;
aud[42621]=16'hd411;
aud[42622]=16'hd421;
aud[42623]=16'hd430;
aud[42624]=16'hd440;
aud[42625]=16'hd450;
aud[42626]=16'hd45f;
aud[42627]=16'hd46f;
aud[42628]=16'hd47f;
aud[42629]=16'hd48f;
aud[42630]=16'hd49e;
aud[42631]=16'hd4ae;
aud[42632]=16'hd4be;
aud[42633]=16'hd4ce;
aud[42634]=16'hd4de;
aud[42635]=16'hd4ed;
aud[42636]=16'hd4fd;
aud[42637]=16'hd50d;
aud[42638]=16'hd51d;
aud[42639]=16'hd52d;
aud[42640]=16'hd53d;
aud[42641]=16'hd54d;
aud[42642]=16'hd55d;
aud[42643]=16'hd56d;
aud[42644]=16'hd57d;
aud[42645]=16'hd58d;
aud[42646]=16'hd59d;
aud[42647]=16'hd5ad;
aud[42648]=16'hd5bd;
aud[42649]=16'hd5cd;
aud[42650]=16'hd5dd;
aud[42651]=16'hd5ee;
aud[42652]=16'hd5fe;
aud[42653]=16'hd60e;
aud[42654]=16'hd61e;
aud[42655]=16'hd62e;
aud[42656]=16'hd63f;
aud[42657]=16'hd64f;
aud[42658]=16'hd65f;
aud[42659]=16'hd66f;
aud[42660]=16'hd680;
aud[42661]=16'hd690;
aud[42662]=16'hd6a0;
aud[42663]=16'hd6b1;
aud[42664]=16'hd6c1;
aud[42665]=16'hd6d2;
aud[42666]=16'hd6e2;
aud[42667]=16'hd6f2;
aud[42668]=16'hd703;
aud[42669]=16'hd713;
aud[42670]=16'hd724;
aud[42671]=16'hd734;
aud[42672]=16'hd745;
aud[42673]=16'hd756;
aud[42674]=16'hd766;
aud[42675]=16'hd777;
aud[42676]=16'hd787;
aud[42677]=16'hd798;
aud[42678]=16'hd7a9;
aud[42679]=16'hd7b9;
aud[42680]=16'hd7ca;
aud[42681]=16'hd7db;
aud[42682]=16'hd7eb;
aud[42683]=16'hd7fc;
aud[42684]=16'hd80d;
aud[42685]=16'hd81e;
aud[42686]=16'hd82e;
aud[42687]=16'hd83f;
aud[42688]=16'hd850;
aud[42689]=16'hd861;
aud[42690]=16'hd872;
aud[42691]=16'hd882;
aud[42692]=16'hd893;
aud[42693]=16'hd8a4;
aud[42694]=16'hd8b5;
aud[42695]=16'hd8c6;
aud[42696]=16'hd8d7;
aud[42697]=16'hd8e8;
aud[42698]=16'hd8f9;
aud[42699]=16'hd90a;
aud[42700]=16'hd91b;
aud[42701]=16'hd92c;
aud[42702]=16'hd93d;
aud[42703]=16'hd94e;
aud[42704]=16'hd95f;
aud[42705]=16'hd970;
aud[42706]=16'hd982;
aud[42707]=16'hd993;
aud[42708]=16'hd9a4;
aud[42709]=16'hd9b5;
aud[42710]=16'hd9c6;
aud[42711]=16'hd9d7;
aud[42712]=16'hd9e9;
aud[42713]=16'hd9fa;
aud[42714]=16'hda0b;
aud[42715]=16'hda1c;
aud[42716]=16'hda2e;
aud[42717]=16'hda3f;
aud[42718]=16'hda50;
aud[42719]=16'hda62;
aud[42720]=16'hda73;
aud[42721]=16'hda84;
aud[42722]=16'hda96;
aud[42723]=16'hdaa7;
aud[42724]=16'hdab9;
aud[42725]=16'hdaca;
aud[42726]=16'hdadc;
aud[42727]=16'hdaed;
aud[42728]=16'hdaff;
aud[42729]=16'hdb10;
aud[42730]=16'hdb22;
aud[42731]=16'hdb33;
aud[42732]=16'hdb45;
aud[42733]=16'hdb56;
aud[42734]=16'hdb68;
aud[42735]=16'hdb79;
aud[42736]=16'hdb8b;
aud[42737]=16'hdb9d;
aud[42738]=16'hdbae;
aud[42739]=16'hdbc0;
aud[42740]=16'hdbd2;
aud[42741]=16'hdbe3;
aud[42742]=16'hdbf5;
aud[42743]=16'hdc07;
aud[42744]=16'hdc19;
aud[42745]=16'hdc2a;
aud[42746]=16'hdc3c;
aud[42747]=16'hdc4e;
aud[42748]=16'hdc60;
aud[42749]=16'hdc72;
aud[42750]=16'hdc83;
aud[42751]=16'hdc95;
aud[42752]=16'hdca7;
aud[42753]=16'hdcb9;
aud[42754]=16'hdccb;
aud[42755]=16'hdcdd;
aud[42756]=16'hdcef;
aud[42757]=16'hdd01;
aud[42758]=16'hdd13;
aud[42759]=16'hdd25;
aud[42760]=16'hdd37;
aud[42761]=16'hdd49;
aud[42762]=16'hdd5b;
aud[42763]=16'hdd6d;
aud[42764]=16'hdd7f;
aud[42765]=16'hdd91;
aud[42766]=16'hdda3;
aud[42767]=16'hddb5;
aud[42768]=16'hddc7;
aud[42769]=16'hddd9;
aud[42770]=16'hddeb;
aud[42771]=16'hddfe;
aud[42772]=16'hde10;
aud[42773]=16'hde22;
aud[42774]=16'hde34;
aud[42775]=16'hde46;
aud[42776]=16'hde59;
aud[42777]=16'hde6b;
aud[42778]=16'hde7d;
aud[42779]=16'hde8f;
aud[42780]=16'hdea2;
aud[42781]=16'hdeb4;
aud[42782]=16'hdec6;
aud[42783]=16'hded9;
aud[42784]=16'hdeeb;
aud[42785]=16'hdefd;
aud[42786]=16'hdf10;
aud[42787]=16'hdf22;
aud[42788]=16'hdf35;
aud[42789]=16'hdf47;
aud[42790]=16'hdf59;
aud[42791]=16'hdf6c;
aud[42792]=16'hdf7e;
aud[42793]=16'hdf91;
aud[42794]=16'hdfa3;
aud[42795]=16'hdfb6;
aud[42796]=16'hdfc8;
aud[42797]=16'hdfdb;
aud[42798]=16'hdfed;
aud[42799]=16'he000;
aud[42800]=16'he013;
aud[42801]=16'he025;
aud[42802]=16'he038;
aud[42803]=16'he04a;
aud[42804]=16'he05d;
aud[42805]=16'he070;
aud[42806]=16'he082;
aud[42807]=16'he095;
aud[42808]=16'he0a8;
aud[42809]=16'he0ba;
aud[42810]=16'he0cd;
aud[42811]=16'he0e0;
aud[42812]=16'he0f3;
aud[42813]=16'he105;
aud[42814]=16'he118;
aud[42815]=16'he12b;
aud[42816]=16'he13e;
aud[42817]=16'he151;
aud[42818]=16'he163;
aud[42819]=16'he176;
aud[42820]=16'he189;
aud[42821]=16'he19c;
aud[42822]=16'he1af;
aud[42823]=16'he1c2;
aud[42824]=16'he1d5;
aud[42825]=16'he1e8;
aud[42826]=16'he1fa;
aud[42827]=16'he20d;
aud[42828]=16'he220;
aud[42829]=16'he233;
aud[42830]=16'he246;
aud[42831]=16'he259;
aud[42832]=16'he26c;
aud[42833]=16'he27f;
aud[42834]=16'he292;
aud[42835]=16'he2a5;
aud[42836]=16'he2b9;
aud[42837]=16'he2cc;
aud[42838]=16'he2df;
aud[42839]=16'he2f2;
aud[42840]=16'he305;
aud[42841]=16'he318;
aud[42842]=16'he32b;
aud[42843]=16'he33e;
aud[42844]=16'he352;
aud[42845]=16'he365;
aud[42846]=16'he378;
aud[42847]=16'he38b;
aud[42848]=16'he39e;
aud[42849]=16'he3b2;
aud[42850]=16'he3c5;
aud[42851]=16'he3d8;
aud[42852]=16'he3eb;
aud[42853]=16'he3ff;
aud[42854]=16'he412;
aud[42855]=16'he425;
aud[42856]=16'he438;
aud[42857]=16'he44c;
aud[42858]=16'he45f;
aud[42859]=16'he473;
aud[42860]=16'he486;
aud[42861]=16'he499;
aud[42862]=16'he4ad;
aud[42863]=16'he4c0;
aud[42864]=16'he4d3;
aud[42865]=16'he4e7;
aud[42866]=16'he4fa;
aud[42867]=16'he50e;
aud[42868]=16'he521;
aud[42869]=16'he535;
aud[42870]=16'he548;
aud[42871]=16'he55c;
aud[42872]=16'he56f;
aud[42873]=16'he583;
aud[42874]=16'he596;
aud[42875]=16'he5aa;
aud[42876]=16'he5bd;
aud[42877]=16'he5d1;
aud[42878]=16'he5e4;
aud[42879]=16'he5f8;
aud[42880]=16'he60c;
aud[42881]=16'he61f;
aud[42882]=16'he633;
aud[42883]=16'he646;
aud[42884]=16'he65a;
aud[42885]=16'he66e;
aud[42886]=16'he681;
aud[42887]=16'he695;
aud[42888]=16'he6a9;
aud[42889]=16'he6bd;
aud[42890]=16'he6d0;
aud[42891]=16'he6e4;
aud[42892]=16'he6f8;
aud[42893]=16'he70b;
aud[42894]=16'he71f;
aud[42895]=16'he733;
aud[42896]=16'he747;
aud[42897]=16'he75b;
aud[42898]=16'he76e;
aud[42899]=16'he782;
aud[42900]=16'he796;
aud[42901]=16'he7aa;
aud[42902]=16'he7be;
aud[42903]=16'he7d1;
aud[42904]=16'he7e5;
aud[42905]=16'he7f9;
aud[42906]=16'he80d;
aud[42907]=16'he821;
aud[42908]=16'he835;
aud[42909]=16'he849;
aud[42910]=16'he85d;
aud[42911]=16'he871;
aud[42912]=16'he885;
aud[42913]=16'he899;
aud[42914]=16'he8ad;
aud[42915]=16'he8c0;
aud[42916]=16'he8d4;
aud[42917]=16'he8e8;
aud[42918]=16'he8fc;
aud[42919]=16'he910;
aud[42920]=16'he925;
aud[42921]=16'he939;
aud[42922]=16'he94d;
aud[42923]=16'he961;
aud[42924]=16'he975;
aud[42925]=16'he989;
aud[42926]=16'he99d;
aud[42927]=16'he9b1;
aud[42928]=16'he9c5;
aud[42929]=16'he9d9;
aud[42930]=16'he9ed;
aud[42931]=16'hea01;
aud[42932]=16'hea16;
aud[42933]=16'hea2a;
aud[42934]=16'hea3e;
aud[42935]=16'hea52;
aud[42936]=16'hea66;
aud[42937]=16'hea7a;
aud[42938]=16'hea8f;
aud[42939]=16'heaa3;
aud[42940]=16'heab7;
aud[42941]=16'heacb;
aud[42942]=16'heae0;
aud[42943]=16'heaf4;
aud[42944]=16'heb08;
aud[42945]=16'heb1c;
aud[42946]=16'heb31;
aud[42947]=16'heb45;
aud[42948]=16'heb59;
aud[42949]=16'heb6e;
aud[42950]=16'heb82;
aud[42951]=16'heb96;
aud[42952]=16'hebab;
aud[42953]=16'hebbf;
aud[42954]=16'hebd3;
aud[42955]=16'hebe8;
aud[42956]=16'hebfc;
aud[42957]=16'hec10;
aud[42958]=16'hec25;
aud[42959]=16'hec39;
aud[42960]=16'hec4d;
aud[42961]=16'hec62;
aud[42962]=16'hec76;
aud[42963]=16'hec8b;
aud[42964]=16'hec9f;
aud[42965]=16'hecb4;
aud[42966]=16'hecc8;
aud[42967]=16'hecdd;
aud[42968]=16'hecf1;
aud[42969]=16'hed05;
aud[42970]=16'hed1a;
aud[42971]=16'hed2e;
aud[42972]=16'hed43;
aud[42973]=16'hed57;
aud[42974]=16'hed6c;
aud[42975]=16'hed81;
aud[42976]=16'hed95;
aud[42977]=16'hedaa;
aud[42978]=16'hedbe;
aud[42979]=16'hedd3;
aud[42980]=16'hede7;
aud[42981]=16'hedfc;
aud[42982]=16'hee10;
aud[42983]=16'hee25;
aud[42984]=16'hee3a;
aud[42985]=16'hee4e;
aud[42986]=16'hee63;
aud[42987]=16'hee77;
aud[42988]=16'hee8c;
aud[42989]=16'heea1;
aud[42990]=16'heeb5;
aud[42991]=16'heeca;
aud[42992]=16'heedf;
aud[42993]=16'heef3;
aud[42994]=16'hef08;
aud[42995]=16'hef1d;
aud[42996]=16'hef31;
aud[42997]=16'hef46;
aud[42998]=16'hef5b;
aud[42999]=16'hef70;
aud[43000]=16'hef84;
aud[43001]=16'hef99;
aud[43002]=16'hefae;
aud[43003]=16'hefc2;
aud[43004]=16'hefd7;
aud[43005]=16'hefec;
aud[43006]=16'hf001;
aud[43007]=16'hf015;
aud[43008]=16'hf02a;
aud[43009]=16'hf03f;
aud[43010]=16'hf054;
aud[43011]=16'hf069;
aud[43012]=16'hf07d;
aud[43013]=16'hf092;
aud[43014]=16'hf0a7;
aud[43015]=16'hf0bc;
aud[43016]=16'hf0d1;
aud[43017]=16'hf0e6;
aud[43018]=16'hf0fa;
aud[43019]=16'hf10f;
aud[43020]=16'hf124;
aud[43021]=16'hf139;
aud[43022]=16'hf14e;
aud[43023]=16'hf163;
aud[43024]=16'hf178;
aud[43025]=16'hf18c;
aud[43026]=16'hf1a1;
aud[43027]=16'hf1b6;
aud[43028]=16'hf1cb;
aud[43029]=16'hf1e0;
aud[43030]=16'hf1f5;
aud[43031]=16'hf20a;
aud[43032]=16'hf21f;
aud[43033]=16'hf234;
aud[43034]=16'hf249;
aud[43035]=16'hf25e;
aud[43036]=16'hf273;
aud[43037]=16'hf288;
aud[43038]=16'hf29d;
aud[43039]=16'hf2b2;
aud[43040]=16'hf2c7;
aud[43041]=16'hf2dc;
aud[43042]=16'hf2f1;
aud[43043]=16'hf306;
aud[43044]=16'hf31b;
aud[43045]=16'hf330;
aud[43046]=16'hf345;
aud[43047]=16'hf35a;
aud[43048]=16'hf36f;
aud[43049]=16'hf384;
aud[43050]=16'hf399;
aud[43051]=16'hf3ae;
aud[43052]=16'hf3c3;
aud[43053]=16'hf3d8;
aud[43054]=16'hf3ed;
aud[43055]=16'hf402;
aud[43056]=16'hf417;
aud[43057]=16'hf42c;
aud[43058]=16'hf441;
aud[43059]=16'hf456;
aud[43060]=16'hf46b;
aud[43061]=16'hf480;
aud[43062]=16'hf496;
aud[43063]=16'hf4ab;
aud[43064]=16'hf4c0;
aud[43065]=16'hf4d5;
aud[43066]=16'hf4ea;
aud[43067]=16'hf4ff;
aud[43068]=16'hf514;
aud[43069]=16'hf529;
aud[43070]=16'hf53f;
aud[43071]=16'hf554;
aud[43072]=16'hf569;
aud[43073]=16'hf57e;
aud[43074]=16'hf593;
aud[43075]=16'hf5a8;
aud[43076]=16'hf5bd;
aud[43077]=16'hf5d3;
aud[43078]=16'hf5e8;
aud[43079]=16'hf5fd;
aud[43080]=16'hf612;
aud[43081]=16'hf627;
aud[43082]=16'hf63d;
aud[43083]=16'hf652;
aud[43084]=16'hf667;
aud[43085]=16'hf67c;
aud[43086]=16'hf691;
aud[43087]=16'hf6a7;
aud[43088]=16'hf6bc;
aud[43089]=16'hf6d1;
aud[43090]=16'hf6e6;
aud[43091]=16'hf6fb;
aud[43092]=16'hf711;
aud[43093]=16'hf726;
aud[43094]=16'hf73b;
aud[43095]=16'hf750;
aud[43096]=16'hf766;
aud[43097]=16'hf77b;
aud[43098]=16'hf790;
aud[43099]=16'hf7a5;
aud[43100]=16'hf7bb;
aud[43101]=16'hf7d0;
aud[43102]=16'hf7e5;
aud[43103]=16'hf7fb;
aud[43104]=16'hf810;
aud[43105]=16'hf825;
aud[43106]=16'hf83a;
aud[43107]=16'hf850;
aud[43108]=16'hf865;
aud[43109]=16'hf87a;
aud[43110]=16'hf890;
aud[43111]=16'hf8a5;
aud[43112]=16'hf8ba;
aud[43113]=16'hf8cf;
aud[43114]=16'hf8e5;
aud[43115]=16'hf8fa;
aud[43116]=16'hf90f;
aud[43117]=16'hf925;
aud[43118]=16'hf93a;
aud[43119]=16'hf94f;
aud[43120]=16'hf965;
aud[43121]=16'hf97a;
aud[43122]=16'hf98f;
aud[43123]=16'hf9a5;
aud[43124]=16'hf9ba;
aud[43125]=16'hf9cf;
aud[43126]=16'hf9e5;
aud[43127]=16'hf9fa;
aud[43128]=16'hfa0f;
aud[43129]=16'hfa25;
aud[43130]=16'hfa3a;
aud[43131]=16'hfa50;
aud[43132]=16'hfa65;
aud[43133]=16'hfa7a;
aud[43134]=16'hfa90;
aud[43135]=16'hfaa5;
aud[43136]=16'hfaba;
aud[43137]=16'hfad0;
aud[43138]=16'hfae5;
aud[43139]=16'hfafb;
aud[43140]=16'hfb10;
aud[43141]=16'hfb25;
aud[43142]=16'hfb3b;
aud[43143]=16'hfb50;
aud[43144]=16'hfb65;
aud[43145]=16'hfb7b;
aud[43146]=16'hfb90;
aud[43147]=16'hfba6;
aud[43148]=16'hfbbb;
aud[43149]=16'hfbd0;
aud[43150]=16'hfbe6;
aud[43151]=16'hfbfb;
aud[43152]=16'hfc11;
aud[43153]=16'hfc26;
aud[43154]=16'hfc3b;
aud[43155]=16'hfc51;
aud[43156]=16'hfc66;
aud[43157]=16'hfc7c;
aud[43158]=16'hfc91;
aud[43159]=16'hfca7;
aud[43160]=16'hfcbc;
aud[43161]=16'hfcd1;
aud[43162]=16'hfce7;
aud[43163]=16'hfcfc;
aud[43164]=16'hfd12;
aud[43165]=16'hfd27;
aud[43166]=16'hfd3c;
aud[43167]=16'hfd52;
aud[43168]=16'hfd67;
aud[43169]=16'hfd7d;
aud[43170]=16'hfd92;
aud[43171]=16'hfda8;
aud[43172]=16'hfdbd;
aud[43173]=16'hfdd2;
aud[43174]=16'hfde8;
aud[43175]=16'hfdfd;
aud[43176]=16'hfe13;
aud[43177]=16'hfe28;
aud[43178]=16'hfe3e;
aud[43179]=16'hfe53;
aud[43180]=16'hfe69;
aud[43181]=16'hfe7e;
aud[43182]=16'hfe93;
aud[43183]=16'hfea9;
aud[43184]=16'hfebe;
aud[43185]=16'hfed4;
aud[43186]=16'hfee9;
aud[43187]=16'hfeff;
aud[43188]=16'hff14;
aud[43189]=16'hff2a;
aud[43190]=16'hff3f;
aud[43191]=16'hff54;
aud[43192]=16'hff6a;
aud[43193]=16'hff7f;
aud[43194]=16'hff95;
aud[43195]=16'hffaa;
aud[43196]=16'hffc0;
aud[43197]=16'hffd5;
aud[43198]=16'hffeb;
aud[43199]=16'h0;
aud[43200]=16'h15;
aud[43201]=16'h2b;
aud[43202]=16'h40;
aud[43203]=16'h56;
aud[43204]=16'h6b;
aud[43205]=16'h81;
aud[43206]=16'h96;
aud[43207]=16'hac;
aud[43208]=16'hc1;
aud[43209]=16'hd6;
aud[43210]=16'hec;
aud[43211]=16'h101;
aud[43212]=16'h117;
aud[43213]=16'h12c;
aud[43214]=16'h142;
aud[43215]=16'h157;
aud[43216]=16'h16d;
aud[43217]=16'h182;
aud[43218]=16'h197;
aud[43219]=16'h1ad;
aud[43220]=16'h1c2;
aud[43221]=16'h1d8;
aud[43222]=16'h1ed;
aud[43223]=16'h203;
aud[43224]=16'h218;
aud[43225]=16'h22e;
aud[43226]=16'h243;
aud[43227]=16'h258;
aud[43228]=16'h26e;
aud[43229]=16'h283;
aud[43230]=16'h299;
aud[43231]=16'h2ae;
aud[43232]=16'h2c4;
aud[43233]=16'h2d9;
aud[43234]=16'h2ee;
aud[43235]=16'h304;
aud[43236]=16'h319;
aud[43237]=16'h32f;
aud[43238]=16'h344;
aud[43239]=16'h359;
aud[43240]=16'h36f;
aud[43241]=16'h384;
aud[43242]=16'h39a;
aud[43243]=16'h3af;
aud[43244]=16'h3c5;
aud[43245]=16'h3da;
aud[43246]=16'h3ef;
aud[43247]=16'h405;
aud[43248]=16'h41a;
aud[43249]=16'h430;
aud[43250]=16'h445;
aud[43251]=16'h45a;
aud[43252]=16'h470;
aud[43253]=16'h485;
aud[43254]=16'h49b;
aud[43255]=16'h4b0;
aud[43256]=16'h4c5;
aud[43257]=16'h4db;
aud[43258]=16'h4f0;
aud[43259]=16'h505;
aud[43260]=16'h51b;
aud[43261]=16'h530;
aud[43262]=16'h546;
aud[43263]=16'h55b;
aud[43264]=16'h570;
aud[43265]=16'h586;
aud[43266]=16'h59b;
aud[43267]=16'h5b0;
aud[43268]=16'h5c6;
aud[43269]=16'h5db;
aud[43270]=16'h5f1;
aud[43271]=16'h606;
aud[43272]=16'h61b;
aud[43273]=16'h631;
aud[43274]=16'h646;
aud[43275]=16'h65b;
aud[43276]=16'h671;
aud[43277]=16'h686;
aud[43278]=16'h69b;
aud[43279]=16'h6b1;
aud[43280]=16'h6c6;
aud[43281]=16'h6db;
aud[43282]=16'h6f1;
aud[43283]=16'h706;
aud[43284]=16'h71b;
aud[43285]=16'h731;
aud[43286]=16'h746;
aud[43287]=16'h75b;
aud[43288]=16'h770;
aud[43289]=16'h786;
aud[43290]=16'h79b;
aud[43291]=16'h7b0;
aud[43292]=16'h7c6;
aud[43293]=16'h7db;
aud[43294]=16'h7f0;
aud[43295]=16'h805;
aud[43296]=16'h81b;
aud[43297]=16'h830;
aud[43298]=16'h845;
aud[43299]=16'h85b;
aud[43300]=16'h870;
aud[43301]=16'h885;
aud[43302]=16'h89a;
aud[43303]=16'h8b0;
aud[43304]=16'h8c5;
aud[43305]=16'h8da;
aud[43306]=16'h8ef;
aud[43307]=16'h905;
aud[43308]=16'h91a;
aud[43309]=16'h92f;
aud[43310]=16'h944;
aud[43311]=16'h959;
aud[43312]=16'h96f;
aud[43313]=16'h984;
aud[43314]=16'h999;
aud[43315]=16'h9ae;
aud[43316]=16'h9c3;
aud[43317]=16'h9d9;
aud[43318]=16'h9ee;
aud[43319]=16'ha03;
aud[43320]=16'ha18;
aud[43321]=16'ha2d;
aud[43322]=16'ha43;
aud[43323]=16'ha58;
aud[43324]=16'ha6d;
aud[43325]=16'ha82;
aud[43326]=16'ha97;
aud[43327]=16'haac;
aud[43328]=16'hac1;
aud[43329]=16'had7;
aud[43330]=16'haec;
aud[43331]=16'hb01;
aud[43332]=16'hb16;
aud[43333]=16'hb2b;
aud[43334]=16'hb40;
aud[43335]=16'hb55;
aud[43336]=16'hb6a;
aud[43337]=16'hb80;
aud[43338]=16'hb95;
aud[43339]=16'hbaa;
aud[43340]=16'hbbf;
aud[43341]=16'hbd4;
aud[43342]=16'hbe9;
aud[43343]=16'hbfe;
aud[43344]=16'hc13;
aud[43345]=16'hc28;
aud[43346]=16'hc3d;
aud[43347]=16'hc52;
aud[43348]=16'hc67;
aud[43349]=16'hc7c;
aud[43350]=16'hc91;
aud[43351]=16'hca6;
aud[43352]=16'hcbb;
aud[43353]=16'hcd0;
aud[43354]=16'hce5;
aud[43355]=16'hcfa;
aud[43356]=16'hd0f;
aud[43357]=16'hd24;
aud[43358]=16'hd39;
aud[43359]=16'hd4e;
aud[43360]=16'hd63;
aud[43361]=16'hd78;
aud[43362]=16'hd8d;
aud[43363]=16'hda2;
aud[43364]=16'hdb7;
aud[43365]=16'hdcc;
aud[43366]=16'hde1;
aud[43367]=16'hdf6;
aud[43368]=16'he0b;
aud[43369]=16'he20;
aud[43370]=16'he35;
aud[43371]=16'he4a;
aud[43372]=16'he5f;
aud[43373]=16'he74;
aud[43374]=16'he88;
aud[43375]=16'he9d;
aud[43376]=16'heb2;
aud[43377]=16'hec7;
aud[43378]=16'hedc;
aud[43379]=16'hef1;
aud[43380]=16'hf06;
aud[43381]=16'hf1a;
aud[43382]=16'hf2f;
aud[43383]=16'hf44;
aud[43384]=16'hf59;
aud[43385]=16'hf6e;
aud[43386]=16'hf83;
aud[43387]=16'hf97;
aud[43388]=16'hfac;
aud[43389]=16'hfc1;
aud[43390]=16'hfd6;
aud[43391]=16'hfeb;
aud[43392]=16'hfff;
aud[43393]=16'h1014;
aud[43394]=16'h1029;
aud[43395]=16'h103e;
aud[43396]=16'h1052;
aud[43397]=16'h1067;
aud[43398]=16'h107c;
aud[43399]=16'h1090;
aud[43400]=16'h10a5;
aud[43401]=16'h10ba;
aud[43402]=16'h10cf;
aud[43403]=16'h10e3;
aud[43404]=16'h10f8;
aud[43405]=16'h110d;
aud[43406]=16'h1121;
aud[43407]=16'h1136;
aud[43408]=16'h114b;
aud[43409]=16'h115f;
aud[43410]=16'h1174;
aud[43411]=16'h1189;
aud[43412]=16'h119d;
aud[43413]=16'h11b2;
aud[43414]=16'h11c6;
aud[43415]=16'h11db;
aud[43416]=16'h11f0;
aud[43417]=16'h1204;
aud[43418]=16'h1219;
aud[43419]=16'h122d;
aud[43420]=16'h1242;
aud[43421]=16'h1256;
aud[43422]=16'h126b;
aud[43423]=16'h127f;
aud[43424]=16'h1294;
aud[43425]=16'h12a9;
aud[43426]=16'h12bd;
aud[43427]=16'h12d2;
aud[43428]=16'h12e6;
aud[43429]=16'h12fb;
aud[43430]=16'h130f;
aud[43431]=16'h1323;
aud[43432]=16'h1338;
aud[43433]=16'h134c;
aud[43434]=16'h1361;
aud[43435]=16'h1375;
aud[43436]=16'h138a;
aud[43437]=16'h139e;
aud[43438]=16'h13b3;
aud[43439]=16'h13c7;
aud[43440]=16'h13db;
aud[43441]=16'h13f0;
aud[43442]=16'h1404;
aud[43443]=16'h1418;
aud[43444]=16'h142d;
aud[43445]=16'h1441;
aud[43446]=16'h1455;
aud[43447]=16'h146a;
aud[43448]=16'h147e;
aud[43449]=16'h1492;
aud[43450]=16'h14a7;
aud[43451]=16'h14bb;
aud[43452]=16'h14cf;
aud[43453]=16'h14e4;
aud[43454]=16'h14f8;
aud[43455]=16'h150c;
aud[43456]=16'h1520;
aud[43457]=16'h1535;
aud[43458]=16'h1549;
aud[43459]=16'h155d;
aud[43460]=16'h1571;
aud[43461]=16'h1586;
aud[43462]=16'h159a;
aud[43463]=16'h15ae;
aud[43464]=16'h15c2;
aud[43465]=16'h15d6;
aud[43466]=16'h15ea;
aud[43467]=16'h15ff;
aud[43468]=16'h1613;
aud[43469]=16'h1627;
aud[43470]=16'h163b;
aud[43471]=16'h164f;
aud[43472]=16'h1663;
aud[43473]=16'h1677;
aud[43474]=16'h168b;
aud[43475]=16'h169f;
aud[43476]=16'h16b3;
aud[43477]=16'h16c7;
aud[43478]=16'h16db;
aud[43479]=16'h16f0;
aud[43480]=16'h1704;
aud[43481]=16'h1718;
aud[43482]=16'h172c;
aud[43483]=16'h1740;
aud[43484]=16'h1753;
aud[43485]=16'h1767;
aud[43486]=16'h177b;
aud[43487]=16'h178f;
aud[43488]=16'h17a3;
aud[43489]=16'h17b7;
aud[43490]=16'h17cb;
aud[43491]=16'h17df;
aud[43492]=16'h17f3;
aud[43493]=16'h1807;
aud[43494]=16'h181b;
aud[43495]=16'h182f;
aud[43496]=16'h1842;
aud[43497]=16'h1856;
aud[43498]=16'h186a;
aud[43499]=16'h187e;
aud[43500]=16'h1892;
aud[43501]=16'h18a5;
aud[43502]=16'h18b9;
aud[43503]=16'h18cd;
aud[43504]=16'h18e1;
aud[43505]=16'h18f5;
aud[43506]=16'h1908;
aud[43507]=16'h191c;
aud[43508]=16'h1930;
aud[43509]=16'h1943;
aud[43510]=16'h1957;
aud[43511]=16'h196b;
aud[43512]=16'h197f;
aud[43513]=16'h1992;
aud[43514]=16'h19a6;
aud[43515]=16'h19ba;
aud[43516]=16'h19cd;
aud[43517]=16'h19e1;
aud[43518]=16'h19f4;
aud[43519]=16'h1a08;
aud[43520]=16'h1a1c;
aud[43521]=16'h1a2f;
aud[43522]=16'h1a43;
aud[43523]=16'h1a56;
aud[43524]=16'h1a6a;
aud[43525]=16'h1a7d;
aud[43526]=16'h1a91;
aud[43527]=16'h1aa4;
aud[43528]=16'h1ab8;
aud[43529]=16'h1acb;
aud[43530]=16'h1adf;
aud[43531]=16'h1af2;
aud[43532]=16'h1b06;
aud[43533]=16'h1b19;
aud[43534]=16'h1b2d;
aud[43535]=16'h1b40;
aud[43536]=16'h1b53;
aud[43537]=16'h1b67;
aud[43538]=16'h1b7a;
aud[43539]=16'h1b8d;
aud[43540]=16'h1ba1;
aud[43541]=16'h1bb4;
aud[43542]=16'h1bc8;
aud[43543]=16'h1bdb;
aud[43544]=16'h1bee;
aud[43545]=16'h1c01;
aud[43546]=16'h1c15;
aud[43547]=16'h1c28;
aud[43548]=16'h1c3b;
aud[43549]=16'h1c4e;
aud[43550]=16'h1c62;
aud[43551]=16'h1c75;
aud[43552]=16'h1c88;
aud[43553]=16'h1c9b;
aud[43554]=16'h1cae;
aud[43555]=16'h1cc2;
aud[43556]=16'h1cd5;
aud[43557]=16'h1ce8;
aud[43558]=16'h1cfb;
aud[43559]=16'h1d0e;
aud[43560]=16'h1d21;
aud[43561]=16'h1d34;
aud[43562]=16'h1d47;
aud[43563]=16'h1d5b;
aud[43564]=16'h1d6e;
aud[43565]=16'h1d81;
aud[43566]=16'h1d94;
aud[43567]=16'h1da7;
aud[43568]=16'h1dba;
aud[43569]=16'h1dcd;
aud[43570]=16'h1de0;
aud[43571]=16'h1df3;
aud[43572]=16'h1e06;
aud[43573]=16'h1e18;
aud[43574]=16'h1e2b;
aud[43575]=16'h1e3e;
aud[43576]=16'h1e51;
aud[43577]=16'h1e64;
aud[43578]=16'h1e77;
aud[43579]=16'h1e8a;
aud[43580]=16'h1e9d;
aud[43581]=16'h1eaf;
aud[43582]=16'h1ec2;
aud[43583]=16'h1ed5;
aud[43584]=16'h1ee8;
aud[43585]=16'h1efb;
aud[43586]=16'h1f0d;
aud[43587]=16'h1f20;
aud[43588]=16'h1f33;
aud[43589]=16'h1f46;
aud[43590]=16'h1f58;
aud[43591]=16'h1f6b;
aud[43592]=16'h1f7e;
aud[43593]=16'h1f90;
aud[43594]=16'h1fa3;
aud[43595]=16'h1fb6;
aud[43596]=16'h1fc8;
aud[43597]=16'h1fdb;
aud[43598]=16'h1fed;
aud[43599]=16'h2000;
aud[43600]=16'h2013;
aud[43601]=16'h2025;
aud[43602]=16'h2038;
aud[43603]=16'h204a;
aud[43604]=16'h205d;
aud[43605]=16'h206f;
aud[43606]=16'h2082;
aud[43607]=16'h2094;
aud[43608]=16'h20a7;
aud[43609]=16'h20b9;
aud[43610]=16'h20cb;
aud[43611]=16'h20de;
aud[43612]=16'h20f0;
aud[43613]=16'h2103;
aud[43614]=16'h2115;
aud[43615]=16'h2127;
aud[43616]=16'h213a;
aud[43617]=16'h214c;
aud[43618]=16'h215e;
aud[43619]=16'h2171;
aud[43620]=16'h2183;
aud[43621]=16'h2195;
aud[43622]=16'h21a7;
aud[43623]=16'h21ba;
aud[43624]=16'h21cc;
aud[43625]=16'h21de;
aud[43626]=16'h21f0;
aud[43627]=16'h2202;
aud[43628]=16'h2215;
aud[43629]=16'h2227;
aud[43630]=16'h2239;
aud[43631]=16'h224b;
aud[43632]=16'h225d;
aud[43633]=16'h226f;
aud[43634]=16'h2281;
aud[43635]=16'h2293;
aud[43636]=16'h22a5;
aud[43637]=16'h22b7;
aud[43638]=16'h22c9;
aud[43639]=16'h22db;
aud[43640]=16'h22ed;
aud[43641]=16'h22ff;
aud[43642]=16'h2311;
aud[43643]=16'h2323;
aud[43644]=16'h2335;
aud[43645]=16'h2347;
aud[43646]=16'h2359;
aud[43647]=16'h236b;
aud[43648]=16'h237d;
aud[43649]=16'h238e;
aud[43650]=16'h23a0;
aud[43651]=16'h23b2;
aud[43652]=16'h23c4;
aud[43653]=16'h23d6;
aud[43654]=16'h23e7;
aud[43655]=16'h23f9;
aud[43656]=16'h240b;
aud[43657]=16'h241d;
aud[43658]=16'h242e;
aud[43659]=16'h2440;
aud[43660]=16'h2452;
aud[43661]=16'h2463;
aud[43662]=16'h2475;
aud[43663]=16'h2487;
aud[43664]=16'h2498;
aud[43665]=16'h24aa;
aud[43666]=16'h24bb;
aud[43667]=16'h24cd;
aud[43668]=16'h24de;
aud[43669]=16'h24f0;
aud[43670]=16'h2501;
aud[43671]=16'h2513;
aud[43672]=16'h2524;
aud[43673]=16'h2536;
aud[43674]=16'h2547;
aud[43675]=16'h2559;
aud[43676]=16'h256a;
aud[43677]=16'h257c;
aud[43678]=16'h258d;
aud[43679]=16'h259e;
aud[43680]=16'h25b0;
aud[43681]=16'h25c1;
aud[43682]=16'h25d2;
aud[43683]=16'h25e4;
aud[43684]=16'h25f5;
aud[43685]=16'h2606;
aud[43686]=16'h2617;
aud[43687]=16'h2629;
aud[43688]=16'h263a;
aud[43689]=16'h264b;
aud[43690]=16'h265c;
aud[43691]=16'h266d;
aud[43692]=16'h267e;
aud[43693]=16'h2690;
aud[43694]=16'h26a1;
aud[43695]=16'h26b2;
aud[43696]=16'h26c3;
aud[43697]=16'h26d4;
aud[43698]=16'h26e5;
aud[43699]=16'h26f6;
aud[43700]=16'h2707;
aud[43701]=16'h2718;
aud[43702]=16'h2729;
aud[43703]=16'h273a;
aud[43704]=16'h274b;
aud[43705]=16'h275c;
aud[43706]=16'h276d;
aud[43707]=16'h277e;
aud[43708]=16'h278e;
aud[43709]=16'h279f;
aud[43710]=16'h27b0;
aud[43711]=16'h27c1;
aud[43712]=16'h27d2;
aud[43713]=16'h27e2;
aud[43714]=16'h27f3;
aud[43715]=16'h2804;
aud[43716]=16'h2815;
aud[43717]=16'h2825;
aud[43718]=16'h2836;
aud[43719]=16'h2847;
aud[43720]=16'h2857;
aud[43721]=16'h2868;
aud[43722]=16'h2879;
aud[43723]=16'h2889;
aud[43724]=16'h289a;
aud[43725]=16'h28aa;
aud[43726]=16'h28bb;
aud[43727]=16'h28cc;
aud[43728]=16'h28dc;
aud[43729]=16'h28ed;
aud[43730]=16'h28fd;
aud[43731]=16'h290e;
aud[43732]=16'h291e;
aud[43733]=16'h292e;
aud[43734]=16'h293f;
aud[43735]=16'h294f;
aud[43736]=16'h2960;
aud[43737]=16'h2970;
aud[43738]=16'h2980;
aud[43739]=16'h2991;
aud[43740]=16'h29a1;
aud[43741]=16'h29b1;
aud[43742]=16'h29c1;
aud[43743]=16'h29d2;
aud[43744]=16'h29e2;
aud[43745]=16'h29f2;
aud[43746]=16'h2a02;
aud[43747]=16'h2a12;
aud[43748]=16'h2a23;
aud[43749]=16'h2a33;
aud[43750]=16'h2a43;
aud[43751]=16'h2a53;
aud[43752]=16'h2a63;
aud[43753]=16'h2a73;
aud[43754]=16'h2a83;
aud[43755]=16'h2a93;
aud[43756]=16'h2aa3;
aud[43757]=16'h2ab3;
aud[43758]=16'h2ac3;
aud[43759]=16'h2ad3;
aud[43760]=16'h2ae3;
aud[43761]=16'h2af3;
aud[43762]=16'h2b03;
aud[43763]=16'h2b13;
aud[43764]=16'h2b22;
aud[43765]=16'h2b32;
aud[43766]=16'h2b42;
aud[43767]=16'h2b52;
aud[43768]=16'h2b62;
aud[43769]=16'h2b71;
aud[43770]=16'h2b81;
aud[43771]=16'h2b91;
aud[43772]=16'h2ba1;
aud[43773]=16'h2bb0;
aud[43774]=16'h2bc0;
aud[43775]=16'h2bd0;
aud[43776]=16'h2bdf;
aud[43777]=16'h2bef;
aud[43778]=16'h2bfe;
aud[43779]=16'h2c0e;
aud[43780]=16'h2c1e;
aud[43781]=16'h2c2d;
aud[43782]=16'h2c3d;
aud[43783]=16'h2c4c;
aud[43784]=16'h2c5c;
aud[43785]=16'h2c6b;
aud[43786]=16'h2c7a;
aud[43787]=16'h2c8a;
aud[43788]=16'h2c99;
aud[43789]=16'h2ca9;
aud[43790]=16'h2cb8;
aud[43791]=16'h2cc7;
aud[43792]=16'h2cd7;
aud[43793]=16'h2ce6;
aud[43794]=16'h2cf5;
aud[43795]=16'h2d04;
aud[43796]=16'h2d14;
aud[43797]=16'h2d23;
aud[43798]=16'h2d32;
aud[43799]=16'h2d41;
aud[43800]=16'h2d50;
aud[43801]=16'h2d60;
aud[43802]=16'h2d6f;
aud[43803]=16'h2d7e;
aud[43804]=16'h2d8d;
aud[43805]=16'h2d9c;
aud[43806]=16'h2dab;
aud[43807]=16'h2dba;
aud[43808]=16'h2dc9;
aud[43809]=16'h2dd8;
aud[43810]=16'h2de7;
aud[43811]=16'h2df6;
aud[43812]=16'h2e05;
aud[43813]=16'h2e14;
aud[43814]=16'h2e22;
aud[43815]=16'h2e31;
aud[43816]=16'h2e40;
aud[43817]=16'h2e4f;
aud[43818]=16'h2e5e;
aud[43819]=16'h2e6d;
aud[43820]=16'h2e7b;
aud[43821]=16'h2e8a;
aud[43822]=16'h2e99;
aud[43823]=16'h2ea7;
aud[43824]=16'h2eb6;
aud[43825]=16'h2ec5;
aud[43826]=16'h2ed3;
aud[43827]=16'h2ee2;
aud[43828]=16'h2ef1;
aud[43829]=16'h2eff;
aud[43830]=16'h2f0e;
aud[43831]=16'h2f1c;
aud[43832]=16'h2f2b;
aud[43833]=16'h2f39;
aud[43834]=16'h2f48;
aud[43835]=16'h2f56;
aud[43836]=16'h2f65;
aud[43837]=16'h2f73;
aud[43838]=16'h2f81;
aud[43839]=16'h2f90;
aud[43840]=16'h2f9e;
aud[43841]=16'h2fac;
aud[43842]=16'h2fbb;
aud[43843]=16'h2fc9;
aud[43844]=16'h2fd7;
aud[43845]=16'h2fe5;
aud[43846]=16'h2ff4;
aud[43847]=16'h3002;
aud[43848]=16'h3010;
aud[43849]=16'h301e;
aud[43850]=16'h302c;
aud[43851]=16'h303a;
aud[43852]=16'h3048;
aud[43853]=16'h3057;
aud[43854]=16'h3065;
aud[43855]=16'h3073;
aud[43856]=16'h3081;
aud[43857]=16'h308f;
aud[43858]=16'h309d;
aud[43859]=16'h30aa;
aud[43860]=16'h30b8;
aud[43861]=16'h30c6;
aud[43862]=16'h30d4;
aud[43863]=16'h30e2;
aud[43864]=16'h30f0;
aud[43865]=16'h30fe;
aud[43866]=16'h310b;
aud[43867]=16'h3119;
aud[43868]=16'h3127;
aud[43869]=16'h3135;
aud[43870]=16'h3142;
aud[43871]=16'h3150;
aud[43872]=16'h315e;
aud[43873]=16'h316b;
aud[43874]=16'h3179;
aud[43875]=16'h3187;
aud[43876]=16'h3194;
aud[43877]=16'h31a2;
aud[43878]=16'h31af;
aud[43879]=16'h31bd;
aud[43880]=16'h31ca;
aud[43881]=16'h31d8;
aud[43882]=16'h31e5;
aud[43883]=16'h31f3;
aud[43884]=16'h3200;
aud[43885]=16'h320d;
aud[43886]=16'h321b;
aud[43887]=16'h3228;
aud[43888]=16'h3235;
aud[43889]=16'h3243;
aud[43890]=16'h3250;
aud[43891]=16'h325d;
aud[43892]=16'h326a;
aud[43893]=16'h3278;
aud[43894]=16'h3285;
aud[43895]=16'h3292;
aud[43896]=16'h329f;
aud[43897]=16'h32ac;
aud[43898]=16'h32b9;
aud[43899]=16'h32c6;
aud[43900]=16'h32d3;
aud[43901]=16'h32e0;
aud[43902]=16'h32ed;
aud[43903]=16'h32fa;
aud[43904]=16'h3307;
aud[43905]=16'h3314;
aud[43906]=16'h3321;
aud[43907]=16'h332e;
aud[43908]=16'h333b;
aud[43909]=16'h3348;
aud[43910]=16'h3355;
aud[43911]=16'h3361;
aud[43912]=16'h336e;
aud[43913]=16'h337b;
aud[43914]=16'h3388;
aud[43915]=16'h3394;
aud[43916]=16'h33a1;
aud[43917]=16'h33ae;
aud[43918]=16'h33ba;
aud[43919]=16'h33c7;
aud[43920]=16'h33d4;
aud[43921]=16'h33e0;
aud[43922]=16'h33ed;
aud[43923]=16'h33f9;
aud[43924]=16'h3406;
aud[43925]=16'h3412;
aud[43926]=16'h341f;
aud[43927]=16'h342b;
aud[43928]=16'h3437;
aud[43929]=16'h3444;
aud[43930]=16'h3450;
aud[43931]=16'h345d;
aud[43932]=16'h3469;
aud[43933]=16'h3475;
aud[43934]=16'h3481;
aud[43935]=16'h348e;
aud[43936]=16'h349a;
aud[43937]=16'h34a6;
aud[43938]=16'h34b2;
aud[43939]=16'h34be;
aud[43940]=16'h34cb;
aud[43941]=16'h34d7;
aud[43942]=16'h34e3;
aud[43943]=16'h34ef;
aud[43944]=16'h34fb;
aud[43945]=16'h3507;
aud[43946]=16'h3513;
aud[43947]=16'h351f;
aud[43948]=16'h352b;
aud[43949]=16'h3537;
aud[43950]=16'h3543;
aud[43951]=16'h354f;
aud[43952]=16'h355a;
aud[43953]=16'h3566;
aud[43954]=16'h3572;
aud[43955]=16'h357e;
aud[43956]=16'h358a;
aud[43957]=16'h3595;
aud[43958]=16'h35a1;
aud[43959]=16'h35ad;
aud[43960]=16'h35b8;
aud[43961]=16'h35c4;
aud[43962]=16'h35d0;
aud[43963]=16'h35db;
aud[43964]=16'h35e7;
aud[43965]=16'h35f2;
aud[43966]=16'h35fe;
aud[43967]=16'h3609;
aud[43968]=16'h3615;
aud[43969]=16'h3620;
aud[43970]=16'h362c;
aud[43971]=16'h3637;
aud[43972]=16'h3643;
aud[43973]=16'h364e;
aud[43974]=16'h3659;
aud[43975]=16'h3665;
aud[43976]=16'h3670;
aud[43977]=16'h367b;
aud[43978]=16'h3686;
aud[43979]=16'h3692;
aud[43980]=16'h369d;
aud[43981]=16'h36a8;
aud[43982]=16'h36b3;
aud[43983]=16'h36be;
aud[43984]=16'h36c9;
aud[43985]=16'h36d4;
aud[43986]=16'h36e0;
aud[43987]=16'h36eb;
aud[43988]=16'h36f6;
aud[43989]=16'h3701;
aud[43990]=16'h370b;
aud[43991]=16'h3716;
aud[43992]=16'h3721;
aud[43993]=16'h372c;
aud[43994]=16'h3737;
aud[43995]=16'h3742;
aud[43996]=16'h374d;
aud[43997]=16'h3757;
aud[43998]=16'h3762;
aud[43999]=16'h376d;
aud[44000]=16'h3778;
aud[44001]=16'h3782;
aud[44002]=16'h378d;
aud[44003]=16'h3798;
aud[44004]=16'h37a2;
aud[44005]=16'h37ad;
aud[44006]=16'h37b7;
aud[44007]=16'h37c2;
aud[44008]=16'h37cc;
aud[44009]=16'h37d7;
aud[44010]=16'h37e1;
aud[44011]=16'h37ec;
aud[44012]=16'h37f6;
aud[44013]=16'h3801;
aud[44014]=16'h380b;
aud[44015]=16'h3815;
aud[44016]=16'h3820;
aud[44017]=16'h382a;
aud[44018]=16'h3834;
aud[44019]=16'h383f;
aud[44020]=16'h3849;
aud[44021]=16'h3853;
aud[44022]=16'h385d;
aud[44023]=16'h3867;
aud[44024]=16'h3871;
aud[44025]=16'h387b;
aud[44026]=16'h3886;
aud[44027]=16'h3890;
aud[44028]=16'h389a;
aud[44029]=16'h38a4;
aud[44030]=16'h38ae;
aud[44031]=16'h38b8;
aud[44032]=16'h38c1;
aud[44033]=16'h38cb;
aud[44034]=16'h38d5;
aud[44035]=16'h38df;
aud[44036]=16'h38e9;
aud[44037]=16'h38f3;
aud[44038]=16'h38fd;
aud[44039]=16'h3906;
aud[44040]=16'h3910;
aud[44041]=16'h391a;
aud[44042]=16'h3923;
aud[44043]=16'h392d;
aud[44044]=16'h3937;
aud[44045]=16'h3940;
aud[44046]=16'h394a;
aud[44047]=16'h3953;
aud[44048]=16'h395d;
aud[44049]=16'h3966;
aud[44050]=16'h3970;
aud[44051]=16'h3979;
aud[44052]=16'h3983;
aud[44053]=16'h398c;
aud[44054]=16'h3995;
aud[44055]=16'h399f;
aud[44056]=16'h39a8;
aud[44057]=16'h39b1;
aud[44058]=16'h39bb;
aud[44059]=16'h39c4;
aud[44060]=16'h39cd;
aud[44061]=16'h39d6;
aud[44062]=16'h39e0;
aud[44063]=16'h39e9;
aud[44064]=16'h39f2;
aud[44065]=16'h39fb;
aud[44066]=16'h3a04;
aud[44067]=16'h3a0d;
aud[44068]=16'h3a16;
aud[44069]=16'h3a1f;
aud[44070]=16'h3a28;
aud[44071]=16'h3a31;
aud[44072]=16'h3a3a;
aud[44073]=16'h3a43;
aud[44074]=16'h3a4c;
aud[44075]=16'h3a54;
aud[44076]=16'h3a5d;
aud[44077]=16'h3a66;
aud[44078]=16'h3a6f;
aud[44079]=16'h3a78;
aud[44080]=16'h3a80;
aud[44081]=16'h3a89;
aud[44082]=16'h3a92;
aud[44083]=16'h3a9a;
aud[44084]=16'h3aa3;
aud[44085]=16'h3aab;
aud[44086]=16'h3ab4;
aud[44087]=16'h3abc;
aud[44088]=16'h3ac5;
aud[44089]=16'h3acd;
aud[44090]=16'h3ad6;
aud[44091]=16'h3ade;
aud[44092]=16'h3ae7;
aud[44093]=16'h3aef;
aud[44094]=16'h3af7;
aud[44095]=16'h3b00;
aud[44096]=16'h3b08;
aud[44097]=16'h3b10;
aud[44098]=16'h3b19;
aud[44099]=16'h3b21;
aud[44100]=16'h3b29;
aud[44101]=16'h3b31;
aud[44102]=16'h3b39;
aud[44103]=16'h3b41;
aud[44104]=16'h3b4a;
aud[44105]=16'h3b52;
aud[44106]=16'h3b5a;
aud[44107]=16'h3b62;
aud[44108]=16'h3b6a;
aud[44109]=16'h3b72;
aud[44110]=16'h3b7a;
aud[44111]=16'h3b81;
aud[44112]=16'h3b89;
aud[44113]=16'h3b91;
aud[44114]=16'h3b99;
aud[44115]=16'h3ba1;
aud[44116]=16'h3ba9;
aud[44117]=16'h3bb0;
aud[44118]=16'h3bb8;
aud[44119]=16'h3bc0;
aud[44120]=16'h3bc7;
aud[44121]=16'h3bcf;
aud[44122]=16'h3bd7;
aud[44123]=16'h3bde;
aud[44124]=16'h3be6;
aud[44125]=16'h3bed;
aud[44126]=16'h3bf5;
aud[44127]=16'h3bfc;
aud[44128]=16'h3c04;
aud[44129]=16'h3c0b;
aud[44130]=16'h3c13;
aud[44131]=16'h3c1a;
aud[44132]=16'h3c21;
aud[44133]=16'h3c29;
aud[44134]=16'h3c30;
aud[44135]=16'h3c37;
aud[44136]=16'h3c3f;
aud[44137]=16'h3c46;
aud[44138]=16'h3c4d;
aud[44139]=16'h3c54;
aud[44140]=16'h3c5b;
aud[44141]=16'h3c63;
aud[44142]=16'h3c6a;
aud[44143]=16'h3c71;
aud[44144]=16'h3c78;
aud[44145]=16'h3c7f;
aud[44146]=16'h3c86;
aud[44147]=16'h3c8d;
aud[44148]=16'h3c94;
aud[44149]=16'h3c9b;
aud[44150]=16'h3ca1;
aud[44151]=16'h3ca8;
aud[44152]=16'h3caf;
aud[44153]=16'h3cb6;
aud[44154]=16'h3cbd;
aud[44155]=16'h3cc3;
aud[44156]=16'h3cca;
aud[44157]=16'h3cd1;
aud[44158]=16'h3cd7;
aud[44159]=16'h3cde;
aud[44160]=16'h3ce5;
aud[44161]=16'h3ceb;
aud[44162]=16'h3cf2;
aud[44163]=16'h3cf8;
aud[44164]=16'h3cff;
aud[44165]=16'h3d05;
aud[44166]=16'h3d0c;
aud[44167]=16'h3d12;
aud[44168]=16'h3d19;
aud[44169]=16'h3d1f;
aud[44170]=16'h3d25;
aud[44171]=16'h3d2c;
aud[44172]=16'h3d32;
aud[44173]=16'h3d38;
aud[44174]=16'h3d3f;
aud[44175]=16'h3d45;
aud[44176]=16'h3d4b;
aud[44177]=16'h3d51;
aud[44178]=16'h3d57;
aud[44179]=16'h3d5d;
aud[44180]=16'h3d63;
aud[44181]=16'h3d69;
aud[44182]=16'h3d6f;
aud[44183]=16'h3d75;
aud[44184]=16'h3d7b;
aud[44185]=16'h3d81;
aud[44186]=16'h3d87;
aud[44187]=16'h3d8d;
aud[44188]=16'h3d93;
aud[44189]=16'h3d99;
aud[44190]=16'h3d9f;
aud[44191]=16'h3da4;
aud[44192]=16'h3daa;
aud[44193]=16'h3db0;
aud[44194]=16'h3db6;
aud[44195]=16'h3dbb;
aud[44196]=16'h3dc1;
aud[44197]=16'h3dc7;
aud[44198]=16'h3dcc;
aud[44199]=16'h3dd2;
aud[44200]=16'h3dd7;
aud[44201]=16'h3ddd;
aud[44202]=16'h3de2;
aud[44203]=16'h3de8;
aud[44204]=16'h3ded;
aud[44205]=16'h3df3;
aud[44206]=16'h3df8;
aud[44207]=16'h3dfd;
aud[44208]=16'h3e03;
aud[44209]=16'h3e08;
aud[44210]=16'h3e0d;
aud[44211]=16'h3e12;
aud[44212]=16'h3e18;
aud[44213]=16'h3e1d;
aud[44214]=16'h3e22;
aud[44215]=16'h3e27;
aud[44216]=16'h3e2c;
aud[44217]=16'h3e31;
aud[44218]=16'h3e36;
aud[44219]=16'h3e3b;
aud[44220]=16'h3e40;
aud[44221]=16'h3e45;
aud[44222]=16'h3e4a;
aud[44223]=16'h3e4f;
aud[44224]=16'h3e54;
aud[44225]=16'h3e59;
aud[44226]=16'h3e5e;
aud[44227]=16'h3e62;
aud[44228]=16'h3e67;
aud[44229]=16'h3e6c;
aud[44230]=16'h3e71;
aud[44231]=16'h3e75;
aud[44232]=16'h3e7a;
aud[44233]=16'h3e7f;
aud[44234]=16'h3e83;
aud[44235]=16'h3e88;
aud[44236]=16'h3e8c;
aud[44237]=16'h3e91;
aud[44238]=16'h3e95;
aud[44239]=16'h3e9a;
aud[44240]=16'h3e9e;
aud[44241]=16'h3ea3;
aud[44242]=16'h3ea7;
aud[44243]=16'h3eac;
aud[44244]=16'h3eb0;
aud[44245]=16'h3eb4;
aud[44246]=16'h3eb9;
aud[44247]=16'h3ebd;
aud[44248]=16'h3ec1;
aud[44249]=16'h3ec5;
aud[44250]=16'h3ec9;
aud[44251]=16'h3ecd;
aud[44252]=16'h3ed2;
aud[44253]=16'h3ed6;
aud[44254]=16'h3eda;
aud[44255]=16'h3ede;
aud[44256]=16'h3ee2;
aud[44257]=16'h3ee6;
aud[44258]=16'h3eea;
aud[44259]=16'h3eee;
aud[44260]=16'h3ef2;
aud[44261]=16'h3ef5;
aud[44262]=16'h3ef9;
aud[44263]=16'h3efd;
aud[44264]=16'h3f01;
aud[44265]=16'h3f05;
aud[44266]=16'h3f08;
aud[44267]=16'h3f0c;
aud[44268]=16'h3f10;
aud[44269]=16'h3f13;
aud[44270]=16'h3f17;
aud[44271]=16'h3f1b;
aud[44272]=16'h3f1e;
aud[44273]=16'h3f22;
aud[44274]=16'h3f25;
aud[44275]=16'h3f29;
aud[44276]=16'h3f2c;
aud[44277]=16'h3f30;
aud[44278]=16'h3f33;
aud[44279]=16'h3f36;
aud[44280]=16'h3f3a;
aud[44281]=16'h3f3d;
aud[44282]=16'h3f40;
aud[44283]=16'h3f43;
aud[44284]=16'h3f47;
aud[44285]=16'h3f4a;
aud[44286]=16'h3f4d;
aud[44287]=16'h3f50;
aud[44288]=16'h3f53;
aud[44289]=16'h3f56;
aud[44290]=16'h3f5a;
aud[44291]=16'h3f5d;
aud[44292]=16'h3f60;
aud[44293]=16'h3f63;
aud[44294]=16'h3f65;
aud[44295]=16'h3f68;
aud[44296]=16'h3f6b;
aud[44297]=16'h3f6e;
aud[44298]=16'h3f71;
aud[44299]=16'h3f74;
aud[44300]=16'h3f77;
aud[44301]=16'h3f79;
aud[44302]=16'h3f7c;
aud[44303]=16'h3f7f;
aud[44304]=16'h3f81;
aud[44305]=16'h3f84;
aud[44306]=16'h3f87;
aud[44307]=16'h3f89;
aud[44308]=16'h3f8c;
aud[44309]=16'h3f8e;
aud[44310]=16'h3f91;
aud[44311]=16'h3f93;
aud[44312]=16'h3f96;
aud[44313]=16'h3f98;
aud[44314]=16'h3f9b;
aud[44315]=16'h3f9d;
aud[44316]=16'h3f9f;
aud[44317]=16'h3fa2;
aud[44318]=16'h3fa4;
aud[44319]=16'h3fa6;
aud[44320]=16'h3fa8;
aud[44321]=16'h3fab;
aud[44322]=16'h3fad;
aud[44323]=16'h3faf;
aud[44324]=16'h3fb1;
aud[44325]=16'h3fb3;
aud[44326]=16'h3fb5;
aud[44327]=16'h3fb7;
aud[44328]=16'h3fb9;
aud[44329]=16'h3fbb;
aud[44330]=16'h3fbd;
aud[44331]=16'h3fbf;
aud[44332]=16'h3fc1;
aud[44333]=16'h3fc3;
aud[44334]=16'h3fc5;
aud[44335]=16'h3fc7;
aud[44336]=16'h3fc8;
aud[44337]=16'h3fca;
aud[44338]=16'h3fcc;
aud[44339]=16'h3fcd;
aud[44340]=16'h3fcf;
aud[44341]=16'h3fd1;
aud[44342]=16'h3fd2;
aud[44343]=16'h3fd4;
aud[44344]=16'h3fd6;
aud[44345]=16'h3fd7;
aud[44346]=16'h3fd9;
aud[44347]=16'h3fda;
aud[44348]=16'h3fdc;
aud[44349]=16'h3fdd;
aud[44350]=16'h3fde;
aud[44351]=16'h3fe0;
aud[44352]=16'h3fe1;
aud[44353]=16'h3fe2;
aud[44354]=16'h3fe4;
aud[44355]=16'h3fe5;
aud[44356]=16'h3fe6;
aud[44357]=16'h3fe7;
aud[44358]=16'h3fe8;
aud[44359]=16'h3fea;
aud[44360]=16'h3feb;
aud[44361]=16'h3fec;
aud[44362]=16'h3fed;
aud[44363]=16'h3fee;
aud[44364]=16'h3fef;
aud[44365]=16'h3ff0;
aud[44366]=16'h3ff1;
aud[44367]=16'h3ff2;
aud[44368]=16'h3ff3;
aud[44369]=16'h3ff3;
aud[44370]=16'h3ff4;
aud[44371]=16'h3ff5;
aud[44372]=16'h3ff6;
aud[44373]=16'h3ff7;
aud[44374]=16'h3ff7;
aud[44375]=16'h3ff8;
aud[44376]=16'h3ff9;
aud[44377]=16'h3ff9;
aud[44378]=16'h3ffa;
aud[44379]=16'h3ffa;
aud[44380]=16'h3ffb;
aud[44381]=16'h3ffb;
aud[44382]=16'h3ffc;
aud[44383]=16'h3ffc;
aud[44384]=16'h3ffd;
aud[44385]=16'h3ffd;
aud[44386]=16'h3ffe;
aud[44387]=16'h3ffe;
aud[44388]=16'h3ffe;
aud[44389]=16'h3fff;
aud[44390]=16'h3fff;
aud[44391]=16'h3fff;
aud[44392]=16'h3fff;
aud[44393]=16'h3fff;
aud[44394]=16'h4000;
aud[44395]=16'h4000;
aud[44396]=16'h4000;
aud[44397]=16'h4000;
aud[44398]=16'h4000;
aud[44399]=16'h4000;
aud[44400]=16'h4000;
aud[44401]=16'h4000;
aud[44402]=16'h4000;
aud[44403]=16'h4000;
aud[44404]=16'h4000;
aud[44405]=16'h3fff;
aud[44406]=16'h3fff;
aud[44407]=16'h3fff;
aud[44408]=16'h3fff;
aud[44409]=16'h3fff;
aud[44410]=16'h3ffe;
aud[44411]=16'h3ffe;
aud[44412]=16'h3ffe;
aud[44413]=16'h3ffd;
aud[44414]=16'h3ffd;
aud[44415]=16'h3ffc;
aud[44416]=16'h3ffc;
aud[44417]=16'h3ffb;
aud[44418]=16'h3ffb;
aud[44419]=16'h3ffa;
aud[44420]=16'h3ffa;
aud[44421]=16'h3ff9;
aud[44422]=16'h3ff9;
aud[44423]=16'h3ff8;
aud[44424]=16'h3ff7;
aud[44425]=16'h3ff7;
aud[44426]=16'h3ff6;
aud[44427]=16'h3ff5;
aud[44428]=16'h3ff4;
aud[44429]=16'h3ff3;
aud[44430]=16'h3ff3;
aud[44431]=16'h3ff2;
aud[44432]=16'h3ff1;
aud[44433]=16'h3ff0;
aud[44434]=16'h3fef;
aud[44435]=16'h3fee;
aud[44436]=16'h3fed;
aud[44437]=16'h3fec;
aud[44438]=16'h3feb;
aud[44439]=16'h3fea;
aud[44440]=16'h3fe8;
aud[44441]=16'h3fe7;
aud[44442]=16'h3fe6;
aud[44443]=16'h3fe5;
aud[44444]=16'h3fe4;
aud[44445]=16'h3fe2;
aud[44446]=16'h3fe1;
aud[44447]=16'h3fe0;
aud[44448]=16'h3fde;
aud[44449]=16'h3fdd;
aud[44450]=16'h3fdc;
aud[44451]=16'h3fda;
aud[44452]=16'h3fd9;
aud[44453]=16'h3fd7;
aud[44454]=16'h3fd6;
aud[44455]=16'h3fd4;
aud[44456]=16'h3fd2;
aud[44457]=16'h3fd1;
aud[44458]=16'h3fcf;
aud[44459]=16'h3fcd;
aud[44460]=16'h3fcc;
aud[44461]=16'h3fca;
aud[44462]=16'h3fc8;
aud[44463]=16'h3fc7;
aud[44464]=16'h3fc5;
aud[44465]=16'h3fc3;
aud[44466]=16'h3fc1;
aud[44467]=16'h3fbf;
aud[44468]=16'h3fbd;
aud[44469]=16'h3fbb;
aud[44470]=16'h3fb9;
aud[44471]=16'h3fb7;
aud[44472]=16'h3fb5;
aud[44473]=16'h3fb3;
aud[44474]=16'h3fb1;
aud[44475]=16'h3faf;
aud[44476]=16'h3fad;
aud[44477]=16'h3fab;
aud[44478]=16'h3fa8;
aud[44479]=16'h3fa6;
aud[44480]=16'h3fa4;
aud[44481]=16'h3fa2;
aud[44482]=16'h3f9f;
aud[44483]=16'h3f9d;
aud[44484]=16'h3f9b;
aud[44485]=16'h3f98;
aud[44486]=16'h3f96;
aud[44487]=16'h3f93;
aud[44488]=16'h3f91;
aud[44489]=16'h3f8e;
aud[44490]=16'h3f8c;
aud[44491]=16'h3f89;
aud[44492]=16'h3f87;
aud[44493]=16'h3f84;
aud[44494]=16'h3f81;
aud[44495]=16'h3f7f;
aud[44496]=16'h3f7c;
aud[44497]=16'h3f79;
aud[44498]=16'h3f77;
aud[44499]=16'h3f74;
aud[44500]=16'h3f71;
aud[44501]=16'h3f6e;
aud[44502]=16'h3f6b;
aud[44503]=16'h3f68;
aud[44504]=16'h3f65;
aud[44505]=16'h3f63;
aud[44506]=16'h3f60;
aud[44507]=16'h3f5d;
aud[44508]=16'h3f5a;
aud[44509]=16'h3f56;
aud[44510]=16'h3f53;
aud[44511]=16'h3f50;
aud[44512]=16'h3f4d;
aud[44513]=16'h3f4a;
aud[44514]=16'h3f47;
aud[44515]=16'h3f43;
aud[44516]=16'h3f40;
aud[44517]=16'h3f3d;
aud[44518]=16'h3f3a;
aud[44519]=16'h3f36;
aud[44520]=16'h3f33;
aud[44521]=16'h3f30;
aud[44522]=16'h3f2c;
aud[44523]=16'h3f29;
aud[44524]=16'h3f25;
aud[44525]=16'h3f22;
aud[44526]=16'h3f1e;
aud[44527]=16'h3f1b;
aud[44528]=16'h3f17;
aud[44529]=16'h3f13;
aud[44530]=16'h3f10;
aud[44531]=16'h3f0c;
aud[44532]=16'h3f08;
aud[44533]=16'h3f05;
aud[44534]=16'h3f01;
aud[44535]=16'h3efd;
aud[44536]=16'h3ef9;
aud[44537]=16'h3ef5;
aud[44538]=16'h3ef2;
aud[44539]=16'h3eee;
aud[44540]=16'h3eea;
aud[44541]=16'h3ee6;
aud[44542]=16'h3ee2;
aud[44543]=16'h3ede;
aud[44544]=16'h3eda;
aud[44545]=16'h3ed6;
aud[44546]=16'h3ed2;
aud[44547]=16'h3ecd;
aud[44548]=16'h3ec9;
aud[44549]=16'h3ec5;
aud[44550]=16'h3ec1;
aud[44551]=16'h3ebd;
aud[44552]=16'h3eb9;
aud[44553]=16'h3eb4;
aud[44554]=16'h3eb0;
aud[44555]=16'h3eac;
aud[44556]=16'h3ea7;
aud[44557]=16'h3ea3;
aud[44558]=16'h3e9e;
aud[44559]=16'h3e9a;
aud[44560]=16'h3e95;
aud[44561]=16'h3e91;
aud[44562]=16'h3e8c;
aud[44563]=16'h3e88;
aud[44564]=16'h3e83;
aud[44565]=16'h3e7f;
aud[44566]=16'h3e7a;
aud[44567]=16'h3e75;
aud[44568]=16'h3e71;
aud[44569]=16'h3e6c;
aud[44570]=16'h3e67;
aud[44571]=16'h3e62;
aud[44572]=16'h3e5e;
aud[44573]=16'h3e59;
aud[44574]=16'h3e54;
aud[44575]=16'h3e4f;
aud[44576]=16'h3e4a;
aud[44577]=16'h3e45;
aud[44578]=16'h3e40;
aud[44579]=16'h3e3b;
aud[44580]=16'h3e36;
aud[44581]=16'h3e31;
aud[44582]=16'h3e2c;
aud[44583]=16'h3e27;
aud[44584]=16'h3e22;
aud[44585]=16'h3e1d;
aud[44586]=16'h3e18;
aud[44587]=16'h3e12;
aud[44588]=16'h3e0d;
aud[44589]=16'h3e08;
aud[44590]=16'h3e03;
aud[44591]=16'h3dfd;
aud[44592]=16'h3df8;
aud[44593]=16'h3df3;
aud[44594]=16'h3ded;
aud[44595]=16'h3de8;
aud[44596]=16'h3de2;
aud[44597]=16'h3ddd;
aud[44598]=16'h3dd7;
aud[44599]=16'h3dd2;
aud[44600]=16'h3dcc;
aud[44601]=16'h3dc7;
aud[44602]=16'h3dc1;
aud[44603]=16'h3dbb;
aud[44604]=16'h3db6;
aud[44605]=16'h3db0;
aud[44606]=16'h3daa;
aud[44607]=16'h3da4;
aud[44608]=16'h3d9f;
aud[44609]=16'h3d99;
aud[44610]=16'h3d93;
aud[44611]=16'h3d8d;
aud[44612]=16'h3d87;
aud[44613]=16'h3d81;
aud[44614]=16'h3d7b;
aud[44615]=16'h3d75;
aud[44616]=16'h3d6f;
aud[44617]=16'h3d69;
aud[44618]=16'h3d63;
aud[44619]=16'h3d5d;
aud[44620]=16'h3d57;
aud[44621]=16'h3d51;
aud[44622]=16'h3d4b;
aud[44623]=16'h3d45;
aud[44624]=16'h3d3f;
aud[44625]=16'h3d38;
aud[44626]=16'h3d32;
aud[44627]=16'h3d2c;
aud[44628]=16'h3d25;
aud[44629]=16'h3d1f;
aud[44630]=16'h3d19;
aud[44631]=16'h3d12;
aud[44632]=16'h3d0c;
aud[44633]=16'h3d05;
aud[44634]=16'h3cff;
aud[44635]=16'h3cf8;
aud[44636]=16'h3cf2;
aud[44637]=16'h3ceb;
aud[44638]=16'h3ce5;
aud[44639]=16'h3cde;
aud[44640]=16'h3cd7;
aud[44641]=16'h3cd1;
aud[44642]=16'h3cca;
aud[44643]=16'h3cc3;
aud[44644]=16'h3cbd;
aud[44645]=16'h3cb6;
aud[44646]=16'h3caf;
aud[44647]=16'h3ca8;
aud[44648]=16'h3ca1;
aud[44649]=16'h3c9b;
aud[44650]=16'h3c94;
aud[44651]=16'h3c8d;
aud[44652]=16'h3c86;
aud[44653]=16'h3c7f;
aud[44654]=16'h3c78;
aud[44655]=16'h3c71;
aud[44656]=16'h3c6a;
aud[44657]=16'h3c63;
aud[44658]=16'h3c5b;
aud[44659]=16'h3c54;
aud[44660]=16'h3c4d;
aud[44661]=16'h3c46;
aud[44662]=16'h3c3f;
aud[44663]=16'h3c37;
aud[44664]=16'h3c30;
aud[44665]=16'h3c29;
aud[44666]=16'h3c21;
aud[44667]=16'h3c1a;
aud[44668]=16'h3c13;
aud[44669]=16'h3c0b;
aud[44670]=16'h3c04;
aud[44671]=16'h3bfc;
aud[44672]=16'h3bf5;
aud[44673]=16'h3bed;
aud[44674]=16'h3be6;
aud[44675]=16'h3bde;
aud[44676]=16'h3bd7;
aud[44677]=16'h3bcf;
aud[44678]=16'h3bc7;
aud[44679]=16'h3bc0;
aud[44680]=16'h3bb8;
aud[44681]=16'h3bb0;
aud[44682]=16'h3ba9;
aud[44683]=16'h3ba1;
aud[44684]=16'h3b99;
aud[44685]=16'h3b91;
aud[44686]=16'h3b89;
aud[44687]=16'h3b81;
aud[44688]=16'h3b7a;
aud[44689]=16'h3b72;
aud[44690]=16'h3b6a;
aud[44691]=16'h3b62;
aud[44692]=16'h3b5a;
aud[44693]=16'h3b52;
aud[44694]=16'h3b4a;
aud[44695]=16'h3b41;
aud[44696]=16'h3b39;
aud[44697]=16'h3b31;
aud[44698]=16'h3b29;
aud[44699]=16'h3b21;
aud[44700]=16'h3b19;
aud[44701]=16'h3b10;
aud[44702]=16'h3b08;
aud[44703]=16'h3b00;
aud[44704]=16'h3af7;
aud[44705]=16'h3aef;
aud[44706]=16'h3ae7;
aud[44707]=16'h3ade;
aud[44708]=16'h3ad6;
aud[44709]=16'h3acd;
aud[44710]=16'h3ac5;
aud[44711]=16'h3abc;
aud[44712]=16'h3ab4;
aud[44713]=16'h3aab;
aud[44714]=16'h3aa3;
aud[44715]=16'h3a9a;
aud[44716]=16'h3a92;
aud[44717]=16'h3a89;
aud[44718]=16'h3a80;
aud[44719]=16'h3a78;
aud[44720]=16'h3a6f;
aud[44721]=16'h3a66;
aud[44722]=16'h3a5d;
aud[44723]=16'h3a54;
aud[44724]=16'h3a4c;
aud[44725]=16'h3a43;
aud[44726]=16'h3a3a;
aud[44727]=16'h3a31;
aud[44728]=16'h3a28;
aud[44729]=16'h3a1f;
aud[44730]=16'h3a16;
aud[44731]=16'h3a0d;
aud[44732]=16'h3a04;
aud[44733]=16'h39fb;
aud[44734]=16'h39f2;
aud[44735]=16'h39e9;
aud[44736]=16'h39e0;
aud[44737]=16'h39d6;
aud[44738]=16'h39cd;
aud[44739]=16'h39c4;
aud[44740]=16'h39bb;
aud[44741]=16'h39b1;
aud[44742]=16'h39a8;
aud[44743]=16'h399f;
aud[44744]=16'h3995;
aud[44745]=16'h398c;
aud[44746]=16'h3983;
aud[44747]=16'h3979;
aud[44748]=16'h3970;
aud[44749]=16'h3966;
aud[44750]=16'h395d;
aud[44751]=16'h3953;
aud[44752]=16'h394a;
aud[44753]=16'h3940;
aud[44754]=16'h3937;
aud[44755]=16'h392d;
aud[44756]=16'h3923;
aud[44757]=16'h391a;
aud[44758]=16'h3910;
aud[44759]=16'h3906;
aud[44760]=16'h38fd;
aud[44761]=16'h38f3;
aud[44762]=16'h38e9;
aud[44763]=16'h38df;
aud[44764]=16'h38d5;
aud[44765]=16'h38cb;
aud[44766]=16'h38c1;
aud[44767]=16'h38b8;
aud[44768]=16'h38ae;
aud[44769]=16'h38a4;
aud[44770]=16'h389a;
aud[44771]=16'h3890;
aud[44772]=16'h3886;
aud[44773]=16'h387b;
aud[44774]=16'h3871;
aud[44775]=16'h3867;
aud[44776]=16'h385d;
aud[44777]=16'h3853;
aud[44778]=16'h3849;
aud[44779]=16'h383f;
aud[44780]=16'h3834;
aud[44781]=16'h382a;
aud[44782]=16'h3820;
aud[44783]=16'h3815;
aud[44784]=16'h380b;
aud[44785]=16'h3801;
aud[44786]=16'h37f6;
aud[44787]=16'h37ec;
aud[44788]=16'h37e1;
aud[44789]=16'h37d7;
aud[44790]=16'h37cc;
aud[44791]=16'h37c2;
aud[44792]=16'h37b7;
aud[44793]=16'h37ad;
aud[44794]=16'h37a2;
aud[44795]=16'h3798;
aud[44796]=16'h378d;
aud[44797]=16'h3782;
aud[44798]=16'h3778;
aud[44799]=16'h376d;
aud[44800]=16'h3762;
aud[44801]=16'h3757;
aud[44802]=16'h374d;
aud[44803]=16'h3742;
aud[44804]=16'h3737;
aud[44805]=16'h372c;
aud[44806]=16'h3721;
aud[44807]=16'h3716;
aud[44808]=16'h370b;
aud[44809]=16'h3701;
aud[44810]=16'h36f6;
aud[44811]=16'h36eb;
aud[44812]=16'h36e0;
aud[44813]=16'h36d4;
aud[44814]=16'h36c9;
aud[44815]=16'h36be;
aud[44816]=16'h36b3;
aud[44817]=16'h36a8;
aud[44818]=16'h369d;
aud[44819]=16'h3692;
aud[44820]=16'h3686;
aud[44821]=16'h367b;
aud[44822]=16'h3670;
aud[44823]=16'h3665;
aud[44824]=16'h3659;
aud[44825]=16'h364e;
aud[44826]=16'h3643;
aud[44827]=16'h3637;
aud[44828]=16'h362c;
aud[44829]=16'h3620;
aud[44830]=16'h3615;
aud[44831]=16'h3609;
aud[44832]=16'h35fe;
aud[44833]=16'h35f2;
aud[44834]=16'h35e7;
aud[44835]=16'h35db;
aud[44836]=16'h35d0;
aud[44837]=16'h35c4;
aud[44838]=16'h35b8;
aud[44839]=16'h35ad;
aud[44840]=16'h35a1;
aud[44841]=16'h3595;
aud[44842]=16'h358a;
aud[44843]=16'h357e;
aud[44844]=16'h3572;
aud[44845]=16'h3566;
aud[44846]=16'h355a;
aud[44847]=16'h354f;
aud[44848]=16'h3543;
aud[44849]=16'h3537;
aud[44850]=16'h352b;
aud[44851]=16'h351f;
aud[44852]=16'h3513;
aud[44853]=16'h3507;
aud[44854]=16'h34fb;
aud[44855]=16'h34ef;
aud[44856]=16'h34e3;
aud[44857]=16'h34d7;
aud[44858]=16'h34cb;
aud[44859]=16'h34be;
aud[44860]=16'h34b2;
aud[44861]=16'h34a6;
aud[44862]=16'h349a;
aud[44863]=16'h348e;
aud[44864]=16'h3481;
aud[44865]=16'h3475;
aud[44866]=16'h3469;
aud[44867]=16'h345d;
aud[44868]=16'h3450;
aud[44869]=16'h3444;
aud[44870]=16'h3437;
aud[44871]=16'h342b;
aud[44872]=16'h341f;
aud[44873]=16'h3412;
aud[44874]=16'h3406;
aud[44875]=16'h33f9;
aud[44876]=16'h33ed;
aud[44877]=16'h33e0;
aud[44878]=16'h33d4;
aud[44879]=16'h33c7;
aud[44880]=16'h33ba;
aud[44881]=16'h33ae;
aud[44882]=16'h33a1;
aud[44883]=16'h3394;
aud[44884]=16'h3388;
aud[44885]=16'h337b;
aud[44886]=16'h336e;
aud[44887]=16'h3361;
aud[44888]=16'h3355;
aud[44889]=16'h3348;
aud[44890]=16'h333b;
aud[44891]=16'h332e;
aud[44892]=16'h3321;
aud[44893]=16'h3314;
aud[44894]=16'h3307;
aud[44895]=16'h32fa;
aud[44896]=16'h32ed;
aud[44897]=16'h32e0;
aud[44898]=16'h32d3;
aud[44899]=16'h32c6;
aud[44900]=16'h32b9;
aud[44901]=16'h32ac;
aud[44902]=16'h329f;
aud[44903]=16'h3292;
aud[44904]=16'h3285;
aud[44905]=16'h3278;
aud[44906]=16'h326a;
aud[44907]=16'h325d;
aud[44908]=16'h3250;
aud[44909]=16'h3243;
aud[44910]=16'h3235;
aud[44911]=16'h3228;
aud[44912]=16'h321b;
aud[44913]=16'h320d;
aud[44914]=16'h3200;
aud[44915]=16'h31f3;
aud[44916]=16'h31e5;
aud[44917]=16'h31d8;
aud[44918]=16'h31ca;
aud[44919]=16'h31bd;
aud[44920]=16'h31af;
aud[44921]=16'h31a2;
aud[44922]=16'h3194;
aud[44923]=16'h3187;
aud[44924]=16'h3179;
aud[44925]=16'h316b;
aud[44926]=16'h315e;
aud[44927]=16'h3150;
aud[44928]=16'h3142;
aud[44929]=16'h3135;
aud[44930]=16'h3127;
aud[44931]=16'h3119;
aud[44932]=16'h310b;
aud[44933]=16'h30fe;
aud[44934]=16'h30f0;
aud[44935]=16'h30e2;
aud[44936]=16'h30d4;
aud[44937]=16'h30c6;
aud[44938]=16'h30b8;
aud[44939]=16'h30aa;
aud[44940]=16'h309d;
aud[44941]=16'h308f;
aud[44942]=16'h3081;
aud[44943]=16'h3073;
aud[44944]=16'h3065;
aud[44945]=16'h3057;
aud[44946]=16'h3048;
aud[44947]=16'h303a;
aud[44948]=16'h302c;
aud[44949]=16'h301e;
aud[44950]=16'h3010;
aud[44951]=16'h3002;
aud[44952]=16'h2ff4;
aud[44953]=16'h2fe5;
aud[44954]=16'h2fd7;
aud[44955]=16'h2fc9;
aud[44956]=16'h2fbb;
aud[44957]=16'h2fac;
aud[44958]=16'h2f9e;
aud[44959]=16'h2f90;
aud[44960]=16'h2f81;
aud[44961]=16'h2f73;
aud[44962]=16'h2f65;
aud[44963]=16'h2f56;
aud[44964]=16'h2f48;
aud[44965]=16'h2f39;
aud[44966]=16'h2f2b;
aud[44967]=16'h2f1c;
aud[44968]=16'h2f0e;
aud[44969]=16'h2eff;
aud[44970]=16'h2ef1;
aud[44971]=16'h2ee2;
aud[44972]=16'h2ed3;
aud[44973]=16'h2ec5;
aud[44974]=16'h2eb6;
aud[44975]=16'h2ea7;
aud[44976]=16'h2e99;
aud[44977]=16'h2e8a;
aud[44978]=16'h2e7b;
aud[44979]=16'h2e6d;
aud[44980]=16'h2e5e;
aud[44981]=16'h2e4f;
aud[44982]=16'h2e40;
aud[44983]=16'h2e31;
aud[44984]=16'h2e22;
aud[44985]=16'h2e14;
aud[44986]=16'h2e05;
aud[44987]=16'h2df6;
aud[44988]=16'h2de7;
aud[44989]=16'h2dd8;
aud[44990]=16'h2dc9;
aud[44991]=16'h2dba;
aud[44992]=16'h2dab;
aud[44993]=16'h2d9c;
aud[44994]=16'h2d8d;
aud[44995]=16'h2d7e;
aud[44996]=16'h2d6f;
aud[44997]=16'h2d60;
aud[44998]=16'h2d50;
aud[44999]=16'h2d41;
aud[45000]=16'h2d32;
aud[45001]=16'h2d23;
aud[45002]=16'h2d14;
aud[45003]=16'h2d04;
aud[45004]=16'h2cf5;
aud[45005]=16'h2ce6;
aud[45006]=16'h2cd7;
aud[45007]=16'h2cc7;
aud[45008]=16'h2cb8;
aud[45009]=16'h2ca9;
aud[45010]=16'h2c99;
aud[45011]=16'h2c8a;
aud[45012]=16'h2c7a;
aud[45013]=16'h2c6b;
aud[45014]=16'h2c5c;
aud[45015]=16'h2c4c;
aud[45016]=16'h2c3d;
aud[45017]=16'h2c2d;
aud[45018]=16'h2c1e;
aud[45019]=16'h2c0e;
aud[45020]=16'h2bfe;
aud[45021]=16'h2bef;
aud[45022]=16'h2bdf;
aud[45023]=16'h2bd0;
aud[45024]=16'h2bc0;
aud[45025]=16'h2bb0;
aud[45026]=16'h2ba1;
aud[45027]=16'h2b91;
aud[45028]=16'h2b81;
aud[45029]=16'h2b71;
aud[45030]=16'h2b62;
aud[45031]=16'h2b52;
aud[45032]=16'h2b42;
aud[45033]=16'h2b32;
aud[45034]=16'h2b22;
aud[45035]=16'h2b13;
aud[45036]=16'h2b03;
aud[45037]=16'h2af3;
aud[45038]=16'h2ae3;
aud[45039]=16'h2ad3;
aud[45040]=16'h2ac3;
aud[45041]=16'h2ab3;
aud[45042]=16'h2aa3;
aud[45043]=16'h2a93;
aud[45044]=16'h2a83;
aud[45045]=16'h2a73;
aud[45046]=16'h2a63;
aud[45047]=16'h2a53;
aud[45048]=16'h2a43;
aud[45049]=16'h2a33;
aud[45050]=16'h2a23;
aud[45051]=16'h2a12;
aud[45052]=16'h2a02;
aud[45053]=16'h29f2;
aud[45054]=16'h29e2;
aud[45055]=16'h29d2;
aud[45056]=16'h29c1;
aud[45057]=16'h29b1;
aud[45058]=16'h29a1;
aud[45059]=16'h2991;
aud[45060]=16'h2980;
aud[45061]=16'h2970;
aud[45062]=16'h2960;
aud[45063]=16'h294f;
aud[45064]=16'h293f;
aud[45065]=16'h292e;
aud[45066]=16'h291e;
aud[45067]=16'h290e;
aud[45068]=16'h28fd;
aud[45069]=16'h28ed;
aud[45070]=16'h28dc;
aud[45071]=16'h28cc;
aud[45072]=16'h28bb;
aud[45073]=16'h28aa;
aud[45074]=16'h289a;
aud[45075]=16'h2889;
aud[45076]=16'h2879;
aud[45077]=16'h2868;
aud[45078]=16'h2857;
aud[45079]=16'h2847;
aud[45080]=16'h2836;
aud[45081]=16'h2825;
aud[45082]=16'h2815;
aud[45083]=16'h2804;
aud[45084]=16'h27f3;
aud[45085]=16'h27e2;
aud[45086]=16'h27d2;
aud[45087]=16'h27c1;
aud[45088]=16'h27b0;
aud[45089]=16'h279f;
aud[45090]=16'h278e;
aud[45091]=16'h277e;
aud[45092]=16'h276d;
aud[45093]=16'h275c;
aud[45094]=16'h274b;
aud[45095]=16'h273a;
aud[45096]=16'h2729;
aud[45097]=16'h2718;
aud[45098]=16'h2707;
aud[45099]=16'h26f6;
aud[45100]=16'h26e5;
aud[45101]=16'h26d4;
aud[45102]=16'h26c3;
aud[45103]=16'h26b2;
aud[45104]=16'h26a1;
aud[45105]=16'h2690;
aud[45106]=16'h267e;
aud[45107]=16'h266d;
aud[45108]=16'h265c;
aud[45109]=16'h264b;
aud[45110]=16'h263a;
aud[45111]=16'h2629;
aud[45112]=16'h2617;
aud[45113]=16'h2606;
aud[45114]=16'h25f5;
aud[45115]=16'h25e4;
aud[45116]=16'h25d2;
aud[45117]=16'h25c1;
aud[45118]=16'h25b0;
aud[45119]=16'h259e;
aud[45120]=16'h258d;
aud[45121]=16'h257c;
aud[45122]=16'h256a;
aud[45123]=16'h2559;
aud[45124]=16'h2547;
aud[45125]=16'h2536;
aud[45126]=16'h2524;
aud[45127]=16'h2513;
aud[45128]=16'h2501;
aud[45129]=16'h24f0;
aud[45130]=16'h24de;
aud[45131]=16'h24cd;
aud[45132]=16'h24bb;
aud[45133]=16'h24aa;
aud[45134]=16'h2498;
aud[45135]=16'h2487;
aud[45136]=16'h2475;
aud[45137]=16'h2463;
aud[45138]=16'h2452;
aud[45139]=16'h2440;
aud[45140]=16'h242e;
aud[45141]=16'h241d;
aud[45142]=16'h240b;
aud[45143]=16'h23f9;
aud[45144]=16'h23e7;
aud[45145]=16'h23d6;
aud[45146]=16'h23c4;
aud[45147]=16'h23b2;
aud[45148]=16'h23a0;
aud[45149]=16'h238e;
aud[45150]=16'h237d;
aud[45151]=16'h236b;
aud[45152]=16'h2359;
aud[45153]=16'h2347;
aud[45154]=16'h2335;
aud[45155]=16'h2323;
aud[45156]=16'h2311;
aud[45157]=16'h22ff;
aud[45158]=16'h22ed;
aud[45159]=16'h22db;
aud[45160]=16'h22c9;
aud[45161]=16'h22b7;
aud[45162]=16'h22a5;
aud[45163]=16'h2293;
aud[45164]=16'h2281;
aud[45165]=16'h226f;
aud[45166]=16'h225d;
aud[45167]=16'h224b;
aud[45168]=16'h2239;
aud[45169]=16'h2227;
aud[45170]=16'h2215;
aud[45171]=16'h2202;
aud[45172]=16'h21f0;
aud[45173]=16'h21de;
aud[45174]=16'h21cc;
aud[45175]=16'h21ba;
aud[45176]=16'h21a7;
aud[45177]=16'h2195;
aud[45178]=16'h2183;
aud[45179]=16'h2171;
aud[45180]=16'h215e;
aud[45181]=16'h214c;
aud[45182]=16'h213a;
aud[45183]=16'h2127;
aud[45184]=16'h2115;
aud[45185]=16'h2103;
aud[45186]=16'h20f0;
aud[45187]=16'h20de;
aud[45188]=16'h20cb;
aud[45189]=16'h20b9;
aud[45190]=16'h20a7;
aud[45191]=16'h2094;
aud[45192]=16'h2082;
aud[45193]=16'h206f;
aud[45194]=16'h205d;
aud[45195]=16'h204a;
aud[45196]=16'h2038;
aud[45197]=16'h2025;
aud[45198]=16'h2013;
aud[45199]=16'h2000;
aud[45200]=16'h1fed;
aud[45201]=16'h1fdb;
aud[45202]=16'h1fc8;
aud[45203]=16'h1fb6;
aud[45204]=16'h1fa3;
aud[45205]=16'h1f90;
aud[45206]=16'h1f7e;
aud[45207]=16'h1f6b;
aud[45208]=16'h1f58;
aud[45209]=16'h1f46;
aud[45210]=16'h1f33;
aud[45211]=16'h1f20;
aud[45212]=16'h1f0d;
aud[45213]=16'h1efb;
aud[45214]=16'h1ee8;
aud[45215]=16'h1ed5;
aud[45216]=16'h1ec2;
aud[45217]=16'h1eaf;
aud[45218]=16'h1e9d;
aud[45219]=16'h1e8a;
aud[45220]=16'h1e77;
aud[45221]=16'h1e64;
aud[45222]=16'h1e51;
aud[45223]=16'h1e3e;
aud[45224]=16'h1e2b;
aud[45225]=16'h1e18;
aud[45226]=16'h1e06;
aud[45227]=16'h1df3;
aud[45228]=16'h1de0;
aud[45229]=16'h1dcd;
aud[45230]=16'h1dba;
aud[45231]=16'h1da7;
aud[45232]=16'h1d94;
aud[45233]=16'h1d81;
aud[45234]=16'h1d6e;
aud[45235]=16'h1d5b;
aud[45236]=16'h1d47;
aud[45237]=16'h1d34;
aud[45238]=16'h1d21;
aud[45239]=16'h1d0e;
aud[45240]=16'h1cfb;
aud[45241]=16'h1ce8;
aud[45242]=16'h1cd5;
aud[45243]=16'h1cc2;
aud[45244]=16'h1cae;
aud[45245]=16'h1c9b;
aud[45246]=16'h1c88;
aud[45247]=16'h1c75;
aud[45248]=16'h1c62;
aud[45249]=16'h1c4e;
aud[45250]=16'h1c3b;
aud[45251]=16'h1c28;
aud[45252]=16'h1c15;
aud[45253]=16'h1c01;
aud[45254]=16'h1bee;
aud[45255]=16'h1bdb;
aud[45256]=16'h1bc8;
aud[45257]=16'h1bb4;
aud[45258]=16'h1ba1;
aud[45259]=16'h1b8d;
aud[45260]=16'h1b7a;
aud[45261]=16'h1b67;
aud[45262]=16'h1b53;
aud[45263]=16'h1b40;
aud[45264]=16'h1b2d;
aud[45265]=16'h1b19;
aud[45266]=16'h1b06;
aud[45267]=16'h1af2;
aud[45268]=16'h1adf;
aud[45269]=16'h1acb;
aud[45270]=16'h1ab8;
aud[45271]=16'h1aa4;
aud[45272]=16'h1a91;
aud[45273]=16'h1a7d;
aud[45274]=16'h1a6a;
aud[45275]=16'h1a56;
aud[45276]=16'h1a43;
aud[45277]=16'h1a2f;
aud[45278]=16'h1a1c;
aud[45279]=16'h1a08;
aud[45280]=16'h19f4;
aud[45281]=16'h19e1;
aud[45282]=16'h19cd;
aud[45283]=16'h19ba;
aud[45284]=16'h19a6;
aud[45285]=16'h1992;
aud[45286]=16'h197f;
aud[45287]=16'h196b;
aud[45288]=16'h1957;
aud[45289]=16'h1943;
aud[45290]=16'h1930;
aud[45291]=16'h191c;
aud[45292]=16'h1908;
aud[45293]=16'h18f5;
aud[45294]=16'h18e1;
aud[45295]=16'h18cd;
aud[45296]=16'h18b9;
aud[45297]=16'h18a5;
aud[45298]=16'h1892;
aud[45299]=16'h187e;
aud[45300]=16'h186a;
aud[45301]=16'h1856;
aud[45302]=16'h1842;
aud[45303]=16'h182f;
aud[45304]=16'h181b;
aud[45305]=16'h1807;
aud[45306]=16'h17f3;
aud[45307]=16'h17df;
aud[45308]=16'h17cb;
aud[45309]=16'h17b7;
aud[45310]=16'h17a3;
aud[45311]=16'h178f;
aud[45312]=16'h177b;
aud[45313]=16'h1767;
aud[45314]=16'h1753;
aud[45315]=16'h1740;
aud[45316]=16'h172c;
aud[45317]=16'h1718;
aud[45318]=16'h1704;
aud[45319]=16'h16f0;
aud[45320]=16'h16db;
aud[45321]=16'h16c7;
aud[45322]=16'h16b3;
aud[45323]=16'h169f;
aud[45324]=16'h168b;
aud[45325]=16'h1677;
aud[45326]=16'h1663;
aud[45327]=16'h164f;
aud[45328]=16'h163b;
aud[45329]=16'h1627;
aud[45330]=16'h1613;
aud[45331]=16'h15ff;
aud[45332]=16'h15ea;
aud[45333]=16'h15d6;
aud[45334]=16'h15c2;
aud[45335]=16'h15ae;
aud[45336]=16'h159a;
aud[45337]=16'h1586;
aud[45338]=16'h1571;
aud[45339]=16'h155d;
aud[45340]=16'h1549;
aud[45341]=16'h1535;
aud[45342]=16'h1520;
aud[45343]=16'h150c;
aud[45344]=16'h14f8;
aud[45345]=16'h14e4;
aud[45346]=16'h14cf;
aud[45347]=16'h14bb;
aud[45348]=16'h14a7;
aud[45349]=16'h1492;
aud[45350]=16'h147e;
aud[45351]=16'h146a;
aud[45352]=16'h1455;
aud[45353]=16'h1441;
aud[45354]=16'h142d;
aud[45355]=16'h1418;
aud[45356]=16'h1404;
aud[45357]=16'h13f0;
aud[45358]=16'h13db;
aud[45359]=16'h13c7;
aud[45360]=16'h13b3;
aud[45361]=16'h139e;
aud[45362]=16'h138a;
aud[45363]=16'h1375;
aud[45364]=16'h1361;
aud[45365]=16'h134c;
aud[45366]=16'h1338;
aud[45367]=16'h1323;
aud[45368]=16'h130f;
aud[45369]=16'h12fb;
aud[45370]=16'h12e6;
aud[45371]=16'h12d2;
aud[45372]=16'h12bd;
aud[45373]=16'h12a9;
aud[45374]=16'h1294;
aud[45375]=16'h127f;
aud[45376]=16'h126b;
aud[45377]=16'h1256;
aud[45378]=16'h1242;
aud[45379]=16'h122d;
aud[45380]=16'h1219;
aud[45381]=16'h1204;
aud[45382]=16'h11f0;
aud[45383]=16'h11db;
aud[45384]=16'h11c6;
aud[45385]=16'h11b2;
aud[45386]=16'h119d;
aud[45387]=16'h1189;
aud[45388]=16'h1174;
aud[45389]=16'h115f;
aud[45390]=16'h114b;
aud[45391]=16'h1136;
aud[45392]=16'h1121;
aud[45393]=16'h110d;
aud[45394]=16'h10f8;
aud[45395]=16'h10e3;
aud[45396]=16'h10cf;
aud[45397]=16'h10ba;
aud[45398]=16'h10a5;
aud[45399]=16'h1090;
aud[45400]=16'h107c;
aud[45401]=16'h1067;
aud[45402]=16'h1052;
aud[45403]=16'h103e;
aud[45404]=16'h1029;
aud[45405]=16'h1014;
aud[45406]=16'hfff;
aud[45407]=16'hfeb;
aud[45408]=16'hfd6;
aud[45409]=16'hfc1;
aud[45410]=16'hfac;
aud[45411]=16'hf97;
aud[45412]=16'hf83;
aud[45413]=16'hf6e;
aud[45414]=16'hf59;
aud[45415]=16'hf44;
aud[45416]=16'hf2f;
aud[45417]=16'hf1a;
aud[45418]=16'hf06;
aud[45419]=16'hef1;
aud[45420]=16'hedc;
aud[45421]=16'hec7;
aud[45422]=16'heb2;
aud[45423]=16'he9d;
aud[45424]=16'he88;
aud[45425]=16'he74;
aud[45426]=16'he5f;
aud[45427]=16'he4a;
aud[45428]=16'he35;
aud[45429]=16'he20;
aud[45430]=16'he0b;
aud[45431]=16'hdf6;
aud[45432]=16'hde1;
aud[45433]=16'hdcc;
aud[45434]=16'hdb7;
aud[45435]=16'hda2;
aud[45436]=16'hd8d;
aud[45437]=16'hd78;
aud[45438]=16'hd63;
aud[45439]=16'hd4e;
aud[45440]=16'hd39;
aud[45441]=16'hd24;
aud[45442]=16'hd0f;
aud[45443]=16'hcfa;
aud[45444]=16'hce5;
aud[45445]=16'hcd0;
aud[45446]=16'hcbb;
aud[45447]=16'hca6;
aud[45448]=16'hc91;
aud[45449]=16'hc7c;
aud[45450]=16'hc67;
aud[45451]=16'hc52;
aud[45452]=16'hc3d;
aud[45453]=16'hc28;
aud[45454]=16'hc13;
aud[45455]=16'hbfe;
aud[45456]=16'hbe9;
aud[45457]=16'hbd4;
aud[45458]=16'hbbf;
aud[45459]=16'hbaa;
aud[45460]=16'hb95;
aud[45461]=16'hb80;
aud[45462]=16'hb6a;
aud[45463]=16'hb55;
aud[45464]=16'hb40;
aud[45465]=16'hb2b;
aud[45466]=16'hb16;
aud[45467]=16'hb01;
aud[45468]=16'haec;
aud[45469]=16'had7;
aud[45470]=16'hac1;
aud[45471]=16'haac;
aud[45472]=16'ha97;
aud[45473]=16'ha82;
aud[45474]=16'ha6d;
aud[45475]=16'ha58;
aud[45476]=16'ha43;
aud[45477]=16'ha2d;
aud[45478]=16'ha18;
aud[45479]=16'ha03;
aud[45480]=16'h9ee;
aud[45481]=16'h9d9;
aud[45482]=16'h9c3;
aud[45483]=16'h9ae;
aud[45484]=16'h999;
aud[45485]=16'h984;
aud[45486]=16'h96f;
aud[45487]=16'h959;
aud[45488]=16'h944;
aud[45489]=16'h92f;
aud[45490]=16'h91a;
aud[45491]=16'h905;
aud[45492]=16'h8ef;
aud[45493]=16'h8da;
aud[45494]=16'h8c5;
aud[45495]=16'h8b0;
aud[45496]=16'h89a;
aud[45497]=16'h885;
aud[45498]=16'h870;
aud[45499]=16'h85b;
aud[45500]=16'h845;
aud[45501]=16'h830;
aud[45502]=16'h81b;
aud[45503]=16'h805;
aud[45504]=16'h7f0;
aud[45505]=16'h7db;
aud[45506]=16'h7c6;
aud[45507]=16'h7b0;
aud[45508]=16'h79b;
aud[45509]=16'h786;
aud[45510]=16'h770;
aud[45511]=16'h75b;
aud[45512]=16'h746;
aud[45513]=16'h731;
aud[45514]=16'h71b;
aud[45515]=16'h706;
aud[45516]=16'h6f1;
aud[45517]=16'h6db;
aud[45518]=16'h6c6;
aud[45519]=16'h6b1;
aud[45520]=16'h69b;
aud[45521]=16'h686;
aud[45522]=16'h671;
aud[45523]=16'h65b;
aud[45524]=16'h646;
aud[45525]=16'h631;
aud[45526]=16'h61b;
aud[45527]=16'h606;
aud[45528]=16'h5f1;
aud[45529]=16'h5db;
aud[45530]=16'h5c6;
aud[45531]=16'h5b0;
aud[45532]=16'h59b;
aud[45533]=16'h586;
aud[45534]=16'h570;
aud[45535]=16'h55b;
aud[45536]=16'h546;
aud[45537]=16'h530;
aud[45538]=16'h51b;
aud[45539]=16'h505;
aud[45540]=16'h4f0;
aud[45541]=16'h4db;
aud[45542]=16'h4c5;
aud[45543]=16'h4b0;
aud[45544]=16'h49b;
aud[45545]=16'h485;
aud[45546]=16'h470;
aud[45547]=16'h45a;
aud[45548]=16'h445;
aud[45549]=16'h430;
aud[45550]=16'h41a;
aud[45551]=16'h405;
aud[45552]=16'h3ef;
aud[45553]=16'h3da;
aud[45554]=16'h3c5;
aud[45555]=16'h3af;
aud[45556]=16'h39a;
aud[45557]=16'h384;
aud[45558]=16'h36f;
aud[45559]=16'h359;
aud[45560]=16'h344;
aud[45561]=16'h32f;
aud[45562]=16'h319;
aud[45563]=16'h304;
aud[45564]=16'h2ee;
aud[45565]=16'h2d9;
aud[45566]=16'h2c4;
aud[45567]=16'h2ae;
aud[45568]=16'h299;
aud[45569]=16'h283;
aud[45570]=16'h26e;
aud[45571]=16'h258;
aud[45572]=16'h243;
aud[45573]=16'h22e;
aud[45574]=16'h218;
aud[45575]=16'h203;
aud[45576]=16'h1ed;
aud[45577]=16'h1d8;
aud[45578]=16'h1c2;
aud[45579]=16'h1ad;
aud[45580]=16'h197;
aud[45581]=16'h182;
aud[45582]=16'h16d;
aud[45583]=16'h157;
aud[45584]=16'h142;
aud[45585]=16'h12c;
aud[45586]=16'h117;
aud[45587]=16'h101;
aud[45588]=16'hec;
aud[45589]=16'hd6;
aud[45590]=16'hc1;
aud[45591]=16'hac;
aud[45592]=16'h96;
aud[45593]=16'h81;
aud[45594]=16'h6b;
aud[45595]=16'h56;
aud[45596]=16'h40;
aud[45597]=16'h2b;
aud[45598]=16'h15;
aud[45599]=16'h0;
aud[45600]=16'hffeb;
aud[45601]=16'hffd5;
aud[45602]=16'hffc0;
aud[45603]=16'hffaa;
aud[45604]=16'hff95;
aud[45605]=16'hff7f;
aud[45606]=16'hff6a;
aud[45607]=16'hff54;
aud[45608]=16'hff3f;
aud[45609]=16'hff2a;
aud[45610]=16'hff14;
aud[45611]=16'hfeff;
aud[45612]=16'hfee9;
aud[45613]=16'hfed4;
aud[45614]=16'hfebe;
aud[45615]=16'hfea9;
aud[45616]=16'hfe93;
aud[45617]=16'hfe7e;
aud[45618]=16'hfe69;
aud[45619]=16'hfe53;
aud[45620]=16'hfe3e;
aud[45621]=16'hfe28;
aud[45622]=16'hfe13;
aud[45623]=16'hfdfd;
aud[45624]=16'hfde8;
aud[45625]=16'hfdd2;
aud[45626]=16'hfdbd;
aud[45627]=16'hfda8;
aud[45628]=16'hfd92;
aud[45629]=16'hfd7d;
aud[45630]=16'hfd67;
aud[45631]=16'hfd52;
aud[45632]=16'hfd3c;
aud[45633]=16'hfd27;
aud[45634]=16'hfd12;
aud[45635]=16'hfcfc;
aud[45636]=16'hfce7;
aud[45637]=16'hfcd1;
aud[45638]=16'hfcbc;
aud[45639]=16'hfca7;
aud[45640]=16'hfc91;
aud[45641]=16'hfc7c;
aud[45642]=16'hfc66;
aud[45643]=16'hfc51;
aud[45644]=16'hfc3b;
aud[45645]=16'hfc26;
aud[45646]=16'hfc11;
aud[45647]=16'hfbfb;
aud[45648]=16'hfbe6;
aud[45649]=16'hfbd0;
aud[45650]=16'hfbbb;
aud[45651]=16'hfba6;
aud[45652]=16'hfb90;
aud[45653]=16'hfb7b;
aud[45654]=16'hfb65;
aud[45655]=16'hfb50;
aud[45656]=16'hfb3b;
aud[45657]=16'hfb25;
aud[45658]=16'hfb10;
aud[45659]=16'hfafb;
aud[45660]=16'hfae5;
aud[45661]=16'hfad0;
aud[45662]=16'hfaba;
aud[45663]=16'hfaa5;
aud[45664]=16'hfa90;
aud[45665]=16'hfa7a;
aud[45666]=16'hfa65;
aud[45667]=16'hfa50;
aud[45668]=16'hfa3a;
aud[45669]=16'hfa25;
aud[45670]=16'hfa0f;
aud[45671]=16'hf9fa;
aud[45672]=16'hf9e5;
aud[45673]=16'hf9cf;
aud[45674]=16'hf9ba;
aud[45675]=16'hf9a5;
aud[45676]=16'hf98f;
aud[45677]=16'hf97a;
aud[45678]=16'hf965;
aud[45679]=16'hf94f;
aud[45680]=16'hf93a;
aud[45681]=16'hf925;
aud[45682]=16'hf90f;
aud[45683]=16'hf8fa;
aud[45684]=16'hf8e5;
aud[45685]=16'hf8cf;
aud[45686]=16'hf8ba;
aud[45687]=16'hf8a5;
aud[45688]=16'hf890;
aud[45689]=16'hf87a;
aud[45690]=16'hf865;
aud[45691]=16'hf850;
aud[45692]=16'hf83a;
aud[45693]=16'hf825;
aud[45694]=16'hf810;
aud[45695]=16'hf7fb;
aud[45696]=16'hf7e5;
aud[45697]=16'hf7d0;
aud[45698]=16'hf7bb;
aud[45699]=16'hf7a5;
aud[45700]=16'hf790;
aud[45701]=16'hf77b;
aud[45702]=16'hf766;
aud[45703]=16'hf750;
aud[45704]=16'hf73b;
aud[45705]=16'hf726;
aud[45706]=16'hf711;
aud[45707]=16'hf6fb;
aud[45708]=16'hf6e6;
aud[45709]=16'hf6d1;
aud[45710]=16'hf6bc;
aud[45711]=16'hf6a7;
aud[45712]=16'hf691;
aud[45713]=16'hf67c;
aud[45714]=16'hf667;
aud[45715]=16'hf652;
aud[45716]=16'hf63d;
aud[45717]=16'hf627;
aud[45718]=16'hf612;
aud[45719]=16'hf5fd;
aud[45720]=16'hf5e8;
aud[45721]=16'hf5d3;
aud[45722]=16'hf5bd;
aud[45723]=16'hf5a8;
aud[45724]=16'hf593;
aud[45725]=16'hf57e;
aud[45726]=16'hf569;
aud[45727]=16'hf554;
aud[45728]=16'hf53f;
aud[45729]=16'hf529;
aud[45730]=16'hf514;
aud[45731]=16'hf4ff;
aud[45732]=16'hf4ea;
aud[45733]=16'hf4d5;
aud[45734]=16'hf4c0;
aud[45735]=16'hf4ab;
aud[45736]=16'hf496;
aud[45737]=16'hf480;
aud[45738]=16'hf46b;
aud[45739]=16'hf456;
aud[45740]=16'hf441;
aud[45741]=16'hf42c;
aud[45742]=16'hf417;
aud[45743]=16'hf402;
aud[45744]=16'hf3ed;
aud[45745]=16'hf3d8;
aud[45746]=16'hf3c3;
aud[45747]=16'hf3ae;
aud[45748]=16'hf399;
aud[45749]=16'hf384;
aud[45750]=16'hf36f;
aud[45751]=16'hf35a;
aud[45752]=16'hf345;
aud[45753]=16'hf330;
aud[45754]=16'hf31b;
aud[45755]=16'hf306;
aud[45756]=16'hf2f1;
aud[45757]=16'hf2dc;
aud[45758]=16'hf2c7;
aud[45759]=16'hf2b2;
aud[45760]=16'hf29d;
aud[45761]=16'hf288;
aud[45762]=16'hf273;
aud[45763]=16'hf25e;
aud[45764]=16'hf249;
aud[45765]=16'hf234;
aud[45766]=16'hf21f;
aud[45767]=16'hf20a;
aud[45768]=16'hf1f5;
aud[45769]=16'hf1e0;
aud[45770]=16'hf1cb;
aud[45771]=16'hf1b6;
aud[45772]=16'hf1a1;
aud[45773]=16'hf18c;
aud[45774]=16'hf178;
aud[45775]=16'hf163;
aud[45776]=16'hf14e;
aud[45777]=16'hf139;
aud[45778]=16'hf124;
aud[45779]=16'hf10f;
aud[45780]=16'hf0fa;
aud[45781]=16'hf0e6;
aud[45782]=16'hf0d1;
aud[45783]=16'hf0bc;
aud[45784]=16'hf0a7;
aud[45785]=16'hf092;
aud[45786]=16'hf07d;
aud[45787]=16'hf069;
aud[45788]=16'hf054;
aud[45789]=16'hf03f;
aud[45790]=16'hf02a;
aud[45791]=16'hf015;
aud[45792]=16'hf001;
aud[45793]=16'hefec;
aud[45794]=16'hefd7;
aud[45795]=16'hefc2;
aud[45796]=16'hefae;
aud[45797]=16'hef99;
aud[45798]=16'hef84;
aud[45799]=16'hef70;
aud[45800]=16'hef5b;
aud[45801]=16'hef46;
aud[45802]=16'hef31;
aud[45803]=16'hef1d;
aud[45804]=16'hef08;
aud[45805]=16'heef3;
aud[45806]=16'heedf;
aud[45807]=16'heeca;
aud[45808]=16'heeb5;
aud[45809]=16'heea1;
aud[45810]=16'hee8c;
aud[45811]=16'hee77;
aud[45812]=16'hee63;
aud[45813]=16'hee4e;
aud[45814]=16'hee3a;
aud[45815]=16'hee25;
aud[45816]=16'hee10;
aud[45817]=16'hedfc;
aud[45818]=16'hede7;
aud[45819]=16'hedd3;
aud[45820]=16'hedbe;
aud[45821]=16'hedaa;
aud[45822]=16'hed95;
aud[45823]=16'hed81;
aud[45824]=16'hed6c;
aud[45825]=16'hed57;
aud[45826]=16'hed43;
aud[45827]=16'hed2e;
aud[45828]=16'hed1a;
aud[45829]=16'hed05;
aud[45830]=16'hecf1;
aud[45831]=16'hecdd;
aud[45832]=16'hecc8;
aud[45833]=16'hecb4;
aud[45834]=16'hec9f;
aud[45835]=16'hec8b;
aud[45836]=16'hec76;
aud[45837]=16'hec62;
aud[45838]=16'hec4d;
aud[45839]=16'hec39;
aud[45840]=16'hec25;
aud[45841]=16'hec10;
aud[45842]=16'hebfc;
aud[45843]=16'hebe8;
aud[45844]=16'hebd3;
aud[45845]=16'hebbf;
aud[45846]=16'hebab;
aud[45847]=16'heb96;
aud[45848]=16'heb82;
aud[45849]=16'heb6e;
aud[45850]=16'heb59;
aud[45851]=16'heb45;
aud[45852]=16'heb31;
aud[45853]=16'heb1c;
aud[45854]=16'heb08;
aud[45855]=16'heaf4;
aud[45856]=16'heae0;
aud[45857]=16'heacb;
aud[45858]=16'heab7;
aud[45859]=16'heaa3;
aud[45860]=16'hea8f;
aud[45861]=16'hea7a;
aud[45862]=16'hea66;
aud[45863]=16'hea52;
aud[45864]=16'hea3e;
aud[45865]=16'hea2a;
aud[45866]=16'hea16;
aud[45867]=16'hea01;
aud[45868]=16'he9ed;
aud[45869]=16'he9d9;
aud[45870]=16'he9c5;
aud[45871]=16'he9b1;
aud[45872]=16'he99d;
aud[45873]=16'he989;
aud[45874]=16'he975;
aud[45875]=16'he961;
aud[45876]=16'he94d;
aud[45877]=16'he939;
aud[45878]=16'he925;
aud[45879]=16'he910;
aud[45880]=16'he8fc;
aud[45881]=16'he8e8;
aud[45882]=16'he8d4;
aud[45883]=16'he8c0;
aud[45884]=16'he8ad;
aud[45885]=16'he899;
aud[45886]=16'he885;
aud[45887]=16'he871;
aud[45888]=16'he85d;
aud[45889]=16'he849;
aud[45890]=16'he835;
aud[45891]=16'he821;
aud[45892]=16'he80d;
aud[45893]=16'he7f9;
aud[45894]=16'he7e5;
aud[45895]=16'he7d1;
aud[45896]=16'he7be;
aud[45897]=16'he7aa;
aud[45898]=16'he796;
aud[45899]=16'he782;
aud[45900]=16'he76e;
aud[45901]=16'he75b;
aud[45902]=16'he747;
aud[45903]=16'he733;
aud[45904]=16'he71f;
aud[45905]=16'he70b;
aud[45906]=16'he6f8;
aud[45907]=16'he6e4;
aud[45908]=16'he6d0;
aud[45909]=16'he6bd;
aud[45910]=16'he6a9;
aud[45911]=16'he695;
aud[45912]=16'he681;
aud[45913]=16'he66e;
aud[45914]=16'he65a;
aud[45915]=16'he646;
aud[45916]=16'he633;
aud[45917]=16'he61f;
aud[45918]=16'he60c;
aud[45919]=16'he5f8;
aud[45920]=16'he5e4;
aud[45921]=16'he5d1;
aud[45922]=16'he5bd;
aud[45923]=16'he5aa;
aud[45924]=16'he596;
aud[45925]=16'he583;
aud[45926]=16'he56f;
aud[45927]=16'he55c;
aud[45928]=16'he548;
aud[45929]=16'he535;
aud[45930]=16'he521;
aud[45931]=16'he50e;
aud[45932]=16'he4fa;
aud[45933]=16'he4e7;
aud[45934]=16'he4d3;
aud[45935]=16'he4c0;
aud[45936]=16'he4ad;
aud[45937]=16'he499;
aud[45938]=16'he486;
aud[45939]=16'he473;
aud[45940]=16'he45f;
aud[45941]=16'he44c;
aud[45942]=16'he438;
aud[45943]=16'he425;
aud[45944]=16'he412;
aud[45945]=16'he3ff;
aud[45946]=16'he3eb;
aud[45947]=16'he3d8;
aud[45948]=16'he3c5;
aud[45949]=16'he3b2;
aud[45950]=16'he39e;
aud[45951]=16'he38b;
aud[45952]=16'he378;
aud[45953]=16'he365;
aud[45954]=16'he352;
aud[45955]=16'he33e;
aud[45956]=16'he32b;
aud[45957]=16'he318;
aud[45958]=16'he305;
aud[45959]=16'he2f2;
aud[45960]=16'he2df;
aud[45961]=16'he2cc;
aud[45962]=16'he2b9;
aud[45963]=16'he2a5;
aud[45964]=16'he292;
aud[45965]=16'he27f;
aud[45966]=16'he26c;
aud[45967]=16'he259;
aud[45968]=16'he246;
aud[45969]=16'he233;
aud[45970]=16'he220;
aud[45971]=16'he20d;
aud[45972]=16'he1fa;
aud[45973]=16'he1e8;
aud[45974]=16'he1d5;
aud[45975]=16'he1c2;
aud[45976]=16'he1af;
aud[45977]=16'he19c;
aud[45978]=16'he189;
aud[45979]=16'he176;
aud[45980]=16'he163;
aud[45981]=16'he151;
aud[45982]=16'he13e;
aud[45983]=16'he12b;
aud[45984]=16'he118;
aud[45985]=16'he105;
aud[45986]=16'he0f3;
aud[45987]=16'he0e0;
aud[45988]=16'he0cd;
aud[45989]=16'he0ba;
aud[45990]=16'he0a8;
aud[45991]=16'he095;
aud[45992]=16'he082;
aud[45993]=16'he070;
aud[45994]=16'he05d;
aud[45995]=16'he04a;
aud[45996]=16'he038;
aud[45997]=16'he025;
aud[45998]=16'he013;
aud[45999]=16'he000;
aud[46000]=16'hdfed;
aud[46001]=16'hdfdb;
aud[46002]=16'hdfc8;
aud[46003]=16'hdfb6;
aud[46004]=16'hdfa3;
aud[46005]=16'hdf91;
aud[46006]=16'hdf7e;
aud[46007]=16'hdf6c;
aud[46008]=16'hdf59;
aud[46009]=16'hdf47;
aud[46010]=16'hdf35;
aud[46011]=16'hdf22;
aud[46012]=16'hdf10;
aud[46013]=16'hdefd;
aud[46014]=16'hdeeb;
aud[46015]=16'hded9;
aud[46016]=16'hdec6;
aud[46017]=16'hdeb4;
aud[46018]=16'hdea2;
aud[46019]=16'hde8f;
aud[46020]=16'hde7d;
aud[46021]=16'hde6b;
aud[46022]=16'hde59;
aud[46023]=16'hde46;
aud[46024]=16'hde34;
aud[46025]=16'hde22;
aud[46026]=16'hde10;
aud[46027]=16'hddfe;
aud[46028]=16'hddeb;
aud[46029]=16'hddd9;
aud[46030]=16'hddc7;
aud[46031]=16'hddb5;
aud[46032]=16'hdda3;
aud[46033]=16'hdd91;
aud[46034]=16'hdd7f;
aud[46035]=16'hdd6d;
aud[46036]=16'hdd5b;
aud[46037]=16'hdd49;
aud[46038]=16'hdd37;
aud[46039]=16'hdd25;
aud[46040]=16'hdd13;
aud[46041]=16'hdd01;
aud[46042]=16'hdcef;
aud[46043]=16'hdcdd;
aud[46044]=16'hdccb;
aud[46045]=16'hdcb9;
aud[46046]=16'hdca7;
aud[46047]=16'hdc95;
aud[46048]=16'hdc83;
aud[46049]=16'hdc72;
aud[46050]=16'hdc60;
aud[46051]=16'hdc4e;
aud[46052]=16'hdc3c;
aud[46053]=16'hdc2a;
aud[46054]=16'hdc19;
aud[46055]=16'hdc07;
aud[46056]=16'hdbf5;
aud[46057]=16'hdbe3;
aud[46058]=16'hdbd2;
aud[46059]=16'hdbc0;
aud[46060]=16'hdbae;
aud[46061]=16'hdb9d;
aud[46062]=16'hdb8b;
aud[46063]=16'hdb79;
aud[46064]=16'hdb68;
aud[46065]=16'hdb56;
aud[46066]=16'hdb45;
aud[46067]=16'hdb33;
aud[46068]=16'hdb22;
aud[46069]=16'hdb10;
aud[46070]=16'hdaff;
aud[46071]=16'hdaed;
aud[46072]=16'hdadc;
aud[46073]=16'hdaca;
aud[46074]=16'hdab9;
aud[46075]=16'hdaa7;
aud[46076]=16'hda96;
aud[46077]=16'hda84;
aud[46078]=16'hda73;
aud[46079]=16'hda62;
aud[46080]=16'hda50;
aud[46081]=16'hda3f;
aud[46082]=16'hda2e;
aud[46083]=16'hda1c;
aud[46084]=16'hda0b;
aud[46085]=16'hd9fa;
aud[46086]=16'hd9e9;
aud[46087]=16'hd9d7;
aud[46088]=16'hd9c6;
aud[46089]=16'hd9b5;
aud[46090]=16'hd9a4;
aud[46091]=16'hd993;
aud[46092]=16'hd982;
aud[46093]=16'hd970;
aud[46094]=16'hd95f;
aud[46095]=16'hd94e;
aud[46096]=16'hd93d;
aud[46097]=16'hd92c;
aud[46098]=16'hd91b;
aud[46099]=16'hd90a;
aud[46100]=16'hd8f9;
aud[46101]=16'hd8e8;
aud[46102]=16'hd8d7;
aud[46103]=16'hd8c6;
aud[46104]=16'hd8b5;
aud[46105]=16'hd8a4;
aud[46106]=16'hd893;
aud[46107]=16'hd882;
aud[46108]=16'hd872;
aud[46109]=16'hd861;
aud[46110]=16'hd850;
aud[46111]=16'hd83f;
aud[46112]=16'hd82e;
aud[46113]=16'hd81e;
aud[46114]=16'hd80d;
aud[46115]=16'hd7fc;
aud[46116]=16'hd7eb;
aud[46117]=16'hd7db;
aud[46118]=16'hd7ca;
aud[46119]=16'hd7b9;
aud[46120]=16'hd7a9;
aud[46121]=16'hd798;
aud[46122]=16'hd787;
aud[46123]=16'hd777;
aud[46124]=16'hd766;
aud[46125]=16'hd756;
aud[46126]=16'hd745;
aud[46127]=16'hd734;
aud[46128]=16'hd724;
aud[46129]=16'hd713;
aud[46130]=16'hd703;
aud[46131]=16'hd6f2;
aud[46132]=16'hd6e2;
aud[46133]=16'hd6d2;
aud[46134]=16'hd6c1;
aud[46135]=16'hd6b1;
aud[46136]=16'hd6a0;
aud[46137]=16'hd690;
aud[46138]=16'hd680;
aud[46139]=16'hd66f;
aud[46140]=16'hd65f;
aud[46141]=16'hd64f;
aud[46142]=16'hd63f;
aud[46143]=16'hd62e;
aud[46144]=16'hd61e;
aud[46145]=16'hd60e;
aud[46146]=16'hd5fe;
aud[46147]=16'hd5ee;
aud[46148]=16'hd5dd;
aud[46149]=16'hd5cd;
aud[46150]=16'hd5bd;
aud[46151]=16'hd5ad;
aud[46152]=16'hd59d;
aud[46153]=16'hd58d;
aud[46154]=16'hd57d;
aud[46155]=16'hd56d;
aud[46156]=16'hd55d;
aud[46157]=16'hd54d;
aud[46158]=16'hd53d;
aud[46159]=16'hd52d;
aud[46160]=16'hd51d;
aud[46161]=16'hd50d;
aud[46162]=16'hd4fd;
aud[46163]=16'hd4ed;
aud[46164]=16'hd4de;
aud[46165]=16'hd4ce;
aud[46166]=16'hd4be;
aud[46167]=16'hd4ae;
aud[46168]=16'hd49e;
aud[46169]=16'hd48f;
aud[46170]=16'hd47f;
aud[46171]=16'hd46f;
aud[46172]=16'hd45f;
aud[46173]=16'hd450;
aud[46174]=16'hd440;
aud[46175]=16'hd430;
aud[46176]=16'hd421;
aud[46177]=16'hd411;
aud[46178]=16'hd402;
aud[46179]=16'hd3f2;
aud[46180]=16'hd3e2;
aud[46181]=16'hd3d3;
aud[46182]=16'hd3c3;
aud[46183]=16'hd3b4;
aud[46184]=16'hd3a4;
aud[46185]=16'hd395;
aud[46186]=16'hd386;
aud[46187]=16'hd376;
aud[46188]=16'hd367;
aud[46189]=16'hd357;
aud[46190]=16'hd348;
aud[46191]=16'hd339;
aud[46192]=16'hd329;
aud[46193]=16'hd31a;
aud[46194]=16'hd30b;
aud[46195]=16'hd2fc;
aud[46196]=16'hd2ec;
aud[46197]=16'hd2dd;
aud[46198]=16'hd2ce;
aud[46199]=16'hd2bf;
aud[46200]=16'hd2b0;
aud[46201]=16'hd2a0;
aud[46202]=16'hd291;
aud[46203]=16'hd282;
aud[46204]=16'hd273;
aud[46205]=16'hd264;
aud[46206]=16'hd255;
aud[46207]=16'hd246;
aud[46208]=16'hd237;
aud[46209]=16'hd228;
aud[46210]=16'hd219;
aud[46211]=16'hd20a;
aud[46212]=16'hd1fb;
aud[46213]=16'hd1ec;
aud[46214]=16'hd1de;
aud[46215]=16'hd1cf;
aud[46216]=16'hd1c0;
aud[46217]=16'hd1b1;
aud[46218]=16'hd1a2;
aud[46219]=16'hd193;
aud[46220]=16'hd185;
aud[46221]=16'hd176;
aud[46222]=16'hd167;
aud[46223]=16'hd159;
aud[46224]=16'hd14a;
aud[46225]=16'hd13b;
aud[46226]=16'hd12d;
aud[46227]=16'hd11e;
aud[46228]=16'hd10f;
aud[46229]=16'hd101;
aud[46230]=16'hd0f2;
aud[46231]=16'hd0e4;
aud[46232]=16'hd0d5;
aud[46233]=16'hd0c7;
aud[46234]=16'hd0b8;
aud[46235]=16'hd0aa;
aud[46236]=16'hd09b;
aud[46237]=16'hd08d;
aud[46238]=16'hd07f;
aud[46239]=16'hd070;
aud[46240]=16'hd062;
aud[46241]=16'hd054;
aud[46242]=16'hd045;
aud[46243]=16'hd037;
aud[46244]=16'hd029;
aud[46245]=16'hd01b;
aud[46246]=16'hd00c;
aud[46247]=16'hcffe;
aud[46248]=16'hcff0;
aud[46249]=16'hcfe2;
aud[46250]=16'hcfd4;
aud[46251]=16'hcfc6;
aud[46252]=16'hcfb8;
aud[46253]=16'hcfa9;
aud[46254]=16'hcf9b;
aud[46255]=16'hcf8d;
aud[46256]=16'hcf7f;
aud[46257]=16'hcf71;
aud[46258]=16'hcf63;
aud[46259]=16'hcf56;
aud[46260]=16'hcf48;
aud[46261]=16'hcf3a;
aud[46262]=16'hcf2c;
aud[46263]=16'hcf1e;
aud[46264]=16'hcf10;
aud[46265]=16'hcf02;
aud[46266]=16'hcef5;
aud[46267]=16'hcee7;
aud[46268]=16'hced9;
aud[46269]=16'hcecb;
aud[46270]=16'hcebe;
aud[46271]=16'hceb0;
aud[46272]=16'hcea2;
aud[46273]=16'hce95;
aud[46274]=16'hce87;
aud[46275]=16'hce79;
aud[46276]=16'hce6c;
aud[46277]=16'hce5e;
aud[46278]=16'hce51;
aud[46279]=16'hce43;
aud[46280]=16'hce36;
aud[46281]=16'hce28;
aud[46282]=16'hce1b;
aud[46283]=16'hce0d;
aud[46284]=16'hce00;
aud[46285]=16'hcdf3;
aud[46286]=16'hcde5;
aud[46287]=16'hcdd8;
aud[46288]=16'hcdcb;
aud[46289]=16'hcdbd;
aud[46290]=16'hcdb0;
aud[46291]=16'hcda3;
aud[46292]=16'hcd96;
aud[46293]=16'hcd88;
aud[46294]=16'hcd7b;
aud[46295]=16'hcd6e;
aud[46296]=16'hcd61;
aud[46297]=16'hcd54;
aud[46298]=16'hcd47;
aud[46299]=16'hcd3a;
aud[46300]=16'hcd2d;
aud[46301]=16'hcd20;
aud[46302]=16'hcd13;
aud[46303]=16'hcd06;
aud[46304]=16'hccf9;
aud[46305]=16'hccec;
aud[46306]=16'hccdf;
aud[46307]=16'hccd2;
aud[46308]=16'hccc5;
aud[46309]=16'hccb8;
aud[46310]=16'hccab;
aud[46311]=16'hcc9f;
aud[46312]=16'hcc92;
aud[46313]=16'hcc85;
aud[46314]=16'hcc78;
aud[46315]=16'hcc6c;
aud[46316]=16'hcc5f;
aud[46317]=16'hcc52;
aud[46318]=16'hcc46;
aud[46319]=16'hcc39;
aud[46320]=16'hcc2c;
aud[46321]=16'hcc20;
aud[46322]=16'hcc13;
aud[46323]=16'hcc07;
aud[46324]=16'hcbfa;
aud[46325]=16'hcbee;
aud[46326]=16'hcbe1;
aud[46327]=16'hcbd5;
aud[46328]=16'hcbc9;
aud[46329]=16'hcbbc;
aud[46330]=16'hcbb0;
aud[46331]=16'hcba3;
aud[46332]=16'hcb97;
aud[46333]=16'hcb8b;
aud[46334]=16'hcb7f;
aud[46335]=16'hcb72;
aud[46336]=16'hcb66;
aud[46337]=16'hcb5a;
aud[46338]=16'hcb4e;
aud[46339]=16'hcb42;
aud[46340]=16'hcb35;
aud[46341]=16'hcb29;
aud[46342]=16'hcb1d;
aud[46343]=16'hcb11;
aud[46344]=16'hcb05;
aud[46345]=16'hcaf9;
aud[46346]=16'hcaed;
aud[46347]=16'hcae1;
aud[46348]=16'hcad5;
aud[46349]=16'hcac9;
aud[46350]=16'hcabd;
aud[46351]=16'hcab1;
aud[46352]=16'hcaa6;
aud[46353]=16'hca9a;
aud[46354]=16'hca8e;
aud[46355]=16'hca82;
aud[46356]=16'hca76;
aud[46357]=16'hca6b;
aud[46358]=16'hca5f;
aud[46359]=16'hca53;
aud[46360]=16'hca48;
aud[46361]=16'hca3c;
aud[46362]=16'hca30;
aud[46363]=16'hca25;
aud[46364]=16'hca19;
aud[46365]=16'hca0e;
aud[46366]=16'hca02;
aud[46367]=16'hc9f7;
aud[46368]=16'hc9eb;
aud[46369]=16'hc9e0;
aud[46370]=16'hc9d4;
aud[46371]=16'hc9c9;
aud[46372]=16'hc9bd;
aud[46373]=16'hc9b2;
aud[46374]=16'hc9a7;
aud[46375]=16'hc99b;
aud[46376]=16'hc990;
aud[46377]=16'hc985;
aud[46378]=16'hc97a;
aud[46379]=16'hc96e;
aud[46380]=16'hc963;
aud[46381]=16'hc958;
aud[46382]=16'hc94d;
aud[46383]=16'hc942;
aud[46384]=16'hc937;
aud[46385]=16'hc92c;
aud[46386]=16'hc920;
aud[46387]=16'hc915;
aud[46388]=16'hc90a;
aud[46389]=16'hc8ff;
aud[46390]=16'hc8f5;
aud[46391]=16'hc8ea;
aud[46392]=16'hc8df;
aud[46393]=16'hc8d4;
aud[46394]=16'hc8c9;
aud[46395]=16'hc8be;
aud[46396]=16'hc8b3;
aud[46397]=16'hc8a9;
aud[46398]=16'hc89e;
aud[46399]=16'hc893;
aud[46400]=16'hc888;
aud[46401]=16'hc87e;
aud[46402]=16'hc873;
aud[46403]=16'hc868;
aud[46404]=16'hc85e;
aud[46405]=16'hc853;
aud[46406]=16'hc849;
aud[46407]=16'hc83e;
aud[46408]=16'hc834;
aud[46409]=16'hc829;
aud[46410]=16'hc81f;
aud[46411]=16'hc814;
aud[46412]=16'hc80a;
aud[46413]=16'hc7ff;
aud[46414]=16'hc7f5;
aud[46415]=16'hc7eb;
aud[46416]=16'hc7e0;
aud[46417]=16'hc7d6;
aud[46418]=16'hc7cc;
aud[46419]=16'hc7c1;
aud[46420]=16'hc7b7;
aud[46421]=16'hc7ad;
aud[46422]=16'hc7a3;
aud[46423]=16'hc799;
aud[46424]=16'hc78f;
aud[46425]=16'hc785;
aud[46426]=16'hc77a;
aud[46427]=16'hc770;
aud[46428]=16'hc766;
aud[46429]=16'hc75c;
aud[46430]=16'hc752;
aud[46431]=16'hc748;
aud[46432]=16'hc73f;
aud[46433]=16'hc735;
aud[46434]=16'hc72b;
aud[46435]=16'hc721;
aud[46436]=16'hc717;
aud[46437]=16'hc70d;
aud[46438]=16'hc703;
aud[46439]=16'hc6fa;
aud[46440]=16'hc6f0;
aud[46441]=16'hc6e6;
aud[46442]=16'hc6dd;
aud[46443]=16'hc6d3;
aud[46444]=16'hc6c9;
aud[46445]=16'hc6c0;
aud[46446]=16'hc6b6;
aud[46447]=16'hc6ad;
aud[46448]=16'hc6a3;
aud[46449]=16'hc69a;
aud[46450]=16'hc690;
aud[46451]=16'hc687;
aud[46452]=16'hc67d;
aud[46453]=16'hc674;
aud[46454]=16'hc66b;
aud[46455]=16'hc661;
aud[46456]=16'hc658;
aud[46457]=16'hc64f;
aud[46458]=16'hc645;
aud[46459]=16'hc63c;
aud[46460]=16'hc633;
aud[46461]=16'hc62a;
aud[46462]=16'hc620;
aud[46463]=16'hc617;
aud[46464]=16'hc60e;
aud[46465]=16'hc605;
aud[46466]=16'hc5fc;
aud[46467]=16'hc5f3;
aud[46468]=16'hc5ea;
aud[46469]=16'hc5e1;
aud[46470]=16'hc5d8;
aud[46471]=16'hc5cf;
aud[46472]=16'hc5c6;
aud[46473]=16'hc5bd;
aud[46474]=16'hc5b4;
aud[46475]=16'hc5ac;
aud[46476]=16'hc5a3;
aud[46477]=16'hc59a;
aud[46478]=16'hc591;
aud[46479]=16'hc588;
aud[46480]=16'hc580;
aud[46481]=16'hc577;
aud[46482]=16'hc56e;
aud[46483]=16'hc566;
aud[46484]=16'hc55d;
aud[46485]=16'hc555;
aud[46486]=16'hc54c;
aud[46487]=16'hc544;
aud[46488]=16'hc53b;
aud[46489]=16'hc533;
aud[46490]=16'hc52a;
aud[46491]=16'hc522;
aud[46492]=16'hc519;
aud[46493]=16'hc511;
aud[46494]=16'hc509;
aud[46495]=16'hc500;
aud[46496]=16'hc4f8;
aud[46497]=16'hc4f0;
aud[46498]=16'hc4e7;
aud[46499]=16'hc4df;
aud[46500]=16'hc4d7;
aud[46501]=16'hc4cf;
aud[46502]=16'hc4c7;
aud[46503]=16'hc4bf;
aud[46504]=16'hc4b6;
aud[46505]=16'hc4ae;
aud[46506]=16'hc4a6;
aud[46507]=16'hc49e;
aud[46508]=16'hc496;
aud[46509]=16'hc48e;
aud[46510]=16'hc486;
aud[46511]=16'hc47f;
aud[46512]=16'hc477;
aud[46513]=16'hc46f;
aud[46514]=16'hc467;
aud[46515]=16'hc45f;
aud[46516]=16'hc457;
aud[46517]=16'hc450;
aud[46518]=16'hc448;
aud[46519]=16'hc440;
aud[46520]=16'hc439;
aud[46521]=16'hc431;
aud[46522]=16'hc429;
aud[46523]=16'hc422;
aud[46524]=16'hc41a;
aud[46525]=16'hc413;
aud[46526]=16'hc40b;
aud[46527]=16'hc404;
aud[46528]=16'hc3fc;
aud[46529]=16'hc3f5;
aud[46530]=16'hc3ed;
aud[46531]=16'hc3e6;
aud[46532]=16'hc3df;
aud[46533]=16'hc3d7;
aud[46534]=16'hc3d0;
aud[46535]=16'hc3c9;
aud[46536]=16'hc3c1;
aud[46537]=16'hc3ba;
aud[46538]=16'hc3b3;
aud[46539]=16'hc3ac;
aud[46540]=16'hc3a5;
aud[46541]=16'hc39d;
aud[46542]=16'hc396;
aud[46543]=16'hc38f;
aud[46544]=16'hc388;
aud[46545]=16'hc381;
aud[46546]=16'hc37a;
aud[46547]=16'hc373;
aud[46548]=16'hc36c;
aud[46549]=16'hc365;
aud[46550]=16'hc35f;
aud[46551]=16'hc358;
aud[46552]=16'hc351;
aud[46553]=16'hc34a;
aud[46554]=16'hc343;
aud[46555]=16'hc33d;
aud[46556]=16'hc336;
aud[46557]=16'hc32f;
aud[46558]=16'hc329;
aud[46559]=16'hc322;
aud[46560]=16'hc31b;
aud[46561]=16'hc315;
aud[46562]=16'hc30e;
aud[46563]=16'hc308;
aud[46564]=16'hc301;
aud[46565]=16'hc2fb;
aud[46566]=16'hc2f4;
aud[46567]=16'hc2ee;
aud[46568]=16'hc2e7;
aud[46569]=16'hc2e1;
aud[46570]=16'hc2db;
aud[46571]=16'hc2d4;
aud[46572]=16'hc2ce;
aud[46573]=16'hc2c8;
aud[46574]=16'hc2c1;
aud[46575]=16'hc2bb;
aud[46576]=16'hc2b5;
aud[46577]=16'hc2af;
aud[46578]=16'hc2a9;
aud[46579]=16'hc2a3;
aud[46580]=16'hc29d;
aud[46581]=16'hc297;
aud[46582]=16'hc291;
aud[46583]=16'hc28b;
aud[46584]=16'hc285;
aud[46585]=16'hc27f;
aud[46586]=16'hc279;
aud[46587]=16'hc273;
aud[46588]=16'hc26d;
aud[46589]=16'hc267;
aud[46590]=16'hc261;
aud[46591]=16'hc25c;
aud[46592]=16'hc256;
aud[46593]=16'hc250;
aud[46594]=16'hc24a;
aud[46595]=16'hc245;
aud[46596]=16'hc23f;
aud[46597]=16'hc239;
aud[46598]=16'hc234;
aud[46599]=16'hc22e;
aud[46600]=16'hc229;
aud[46601]=16'hc223;
aud[46602]=16'hc21e;
aud[46603]=16'hc218;
aud[46604]=16'hc213;
aud[46605]=16'hc20d;
aud[46606]=16'hc208;
aud[46607]=16'hc203;
aud[46608]=16'hc1fd;
aud[46609]=16'hc1f8;
aud[46610]=16'hc1f3;
aud[46611]=16'hc1ee;
aud[46612]=16'hc1e8;
aud[46613]=16'hc1e3;
aud[46614]=16'hc1de;
aud[46615]=16'hc1d9;
aud[46616]=16'hc1d4;
aud[46617]=16'hc1cf;
aud[46618]=16'hc1ca;
aud[46619]=16'hc1c5;
aud[46620]=16'hc1c0;
aud[46621]=16'hc1bb;
aud[46622]=16'hc1b6;
aud[46623]=16'hc1b1;
aud[46624]=16'hc1ac;
aud[46625]=16'hc1a7;
aud[46626]=16'hc1a2;
aud[46627]=16'hc19e;
aud[46628]=16'hc199;
aud[46629]=16'hc194;
aud[46630]=16'hc18f;
aud[46631]=16'hc18b;
aud[46632]=16'hc186;
aud[46633]=16'hc181;
aud[46634]=16'hc17d;
aud[46635]=16'hc178;
aud[46636]=16'hc174;
aud[46637]=16'hc16f;
aud[46638]=16'hc16b;
aud[46639]=16'hc166;
aud[46640]=16'hc162;
aud[46641]=16'hc15d;
aud[46642]=16'hc159;
aud[46643]=16'hc154;
aud[46644]=16'hc150;
aud[46645]=16'hc14c;
aud[46646]=16'hc147;
aud[46647]=16'hc143;
aud[46648]=16'hc13f;
aud[46649]=16'hc13b;
aud[46650]=16'hc137;
aud[46651]=16'hc133;
aud[46652]=16'hc12e;
aud[46653]=16'hc12a;
aud[46654]=16'hc126;
aud[46655]=16'hc122;
aud[46656]=16'hc11e;
aud[46657]=16'hc11a;
aud[46658]=16'hc116;
aud[46659]=16'hc112;
aud[46660]=16'hc10e;
aud[46661]=16'hc10b;
aud[46662]=16'hc107;
aud[46663]=16'hc103;
aud[46664]=16'hc0ff;
aud[46665]=16'hc0fb;
aud[46666]=16'hc0f8;
aud[46667]=16'hc0f4;
aud[46668]=16'hc0f0;
aud[46669]=16'hc0ed;
aud[46670]=16'hc0e9;
aud[46671]=16'hc0e5;
aud[46672]=16'hc0e2;
aud[46673]=16'hc0de;
aud[46674]=16'hc0db;
aud[46675]=16'hc0d7;
aud[46676]=16'hc0d4;
aud[46677]=16'hc0d0;
aud[46678]=16'hc0cd;
aud[46679]=16'hc0ca;
aud[46680]=16'hc0c6;
aud[46681]=16'hc0c3;
aud[46682]=16'hc0c0;
aud[46683]=16'hc0bd;
aud[46684]=16'hc0b9;
aud[46685]=16'hc0b6;
aud[46686]=16'hc0b3;
aud[46687]=16'hc0b0;
aud[46688]=16'hc0ad;
aud[46689]=16'hc0aa;
aud[46690]=16'hc0a6;
aud[46691]=16'hc0a3;
aud[46692]=16'hc0a0;
aud[46693]=16'hc09d;
aud[46694]=16'hc09b;
aud[46695]=16'hc098;
aud[46696]=16'hc095;
aud[46697]=16'hc092;
aud[46698]=16'hc08f;
aud[46699]=16'hc08c;
aud[46700]=16'hc089;
aud[46701]=16'hc087;
aud[46702]=16'hc084;
aud[46703]=16'hc081;
aud[46704]=16'hc07f;
aud[46705]=16'hc07c;
aud[46706]=16'hc079;
aud[46707]=16'hc077;
aud[46708]=16'hc074;
aud[46709]=16'hc072;
aud[46710]=16'hc06f;
aud[46711]=16'hc06d;
aud[46712]=16'hc06a;
aud[46713]=16'hc068;
aud[46714]=16'hc065;
aud[46715]=16'hc063;
aud[46716]=16'hc061;
aud[46717]=16'hc05e;
aud[46718]=16'hc05c;
aud[46719]=16'hc05a;
aud[46720]=16'hc058;
aud[46721]=16'hc055;
aud[46722]=16'hc053;
aud[46723]=16'hc051;
aud[46724]=16'hc04f;
aud[46725]=16'hc04d;
aud[46726]=16'hc04b;
aud[46727]=16'hc049;
aud[46728]=16'hc047;
aud[46729]=16'hc045;
aud[46730]=16'hc043;
aud[46731]=16'hc041;
aud[46732]=16'hc03f;
aud[46733]=16'hc03d;
aud[46734]=16'hc03b;
aud[46735]=16'hc039;
aud[46736]=16'hc038;
aud[46737]=16'hc036;
aud[46738]=16'hc034;
aud[46739]=16'hc033;
aud[46740]=16'hc031;
aud[46741]=16'hc02f;
aud[46742]=16'hc02e;
aud[46743]=16'hc02c;
aud[46744]=16'hc02a;
aud[46745]=16'hc029;
aud[46746]=16'hc027;
aud[46747]=16'hc026;
aud[46748]=16'hc024;
aud[46749]=16'hc023;
aud[46750]=16'hc022;
aud[46751]=16'hc020;
aud[46752]=16'hc01f;
aud[46753]=16'hc01e;
aud[46754]=16'hc01c;
aud[46755]=16'hc01b;
aud[46756]=16'hc01a;
aud[46757]=16'hc019;
aud[46758]=16'hc018;
aud[46759]=16'hc016;
aud[46760]=16'hc015;
aud[46761]=16'hc014;
aud[46762]=16'hc013;
aud[46763]=16'hc012;
aud[46764]=16'hc011;
aud[46765]=16'hc010;
aud[46766]=16'hc00f;
aud[46767]=16'hc00e;
aud[46768]=16'hc00d;
aud[46769]=16'hc00d;
aud[46770]=16'hc00c;
aud[46771]=16'hc00b;
aud[46772]=16'hc00a;
aud[46773]=16'hc009;
aud[46774]=16'hc009;
aud[46775]=16'hc008;
aud[46776]=16'hc007;
aud[46777]=16'hc007;
aud[46778]=16'hc006;
aud[46779]=16'hc006;
aud[46780]=16'hc005;
aud[46781]=16'hc005;
aud[46782]=16'hc004;
aud[46783]=16'hc004;
aud[46784]=16'hc003;
aud[46785]=16'hc003;
aud[46786]=16'hc002;
aud[46787]=16'hc002;
aud[46788]=16'hc002;
aud[46789]=16'hc001;
aud[46790]=16'hc001;
aud[46791]=16'hc001;
aud[46792]=16'hc001;
aud[46793]=16'hc001;
aud[46794]=16'hc000;
aud[46795]=16'hc000;
aud[46796]=16'hc000;
aud[46797]=16'hc000;
aud[46798]=16'hc000;
aud[46799]=16'hc000;
aud[46800]=16'hc000;
aud[46801]=16'hc000;
aud[46802]=16'hc000;
aud[46803]=16'hc000;
aud[46804]=16'hc000;
aud[46805]=16'hc001;
aud[46806]=16'hc001;
aud[46807]=16'hc001;
aud[46808]=16'hc001;
aud[46809]=16'hc001;
aud[46810]=16'hc002;
aud[46811]=16'hc002;
aud[46812]=16'hc002;
aud[46813]=16'hc003;
aud[46814]=16'hc003;
aud[46815]=16'hc004;
aud[46816]=16'hc004;
aud[46817]=16'hc005;
aud[46818]=16'hc005;
aud[46819]=16'hc006;
aud[46820]=16'hc006;
aud[46821]=16'hc007;
aud[46822]=16'hc007;
aud[46823]=16'hc008;
aud[46824]=16'hc009;
aud[46825]=16'hc009;
aud[46826]=16'hc00a;
aud[46827]=16'hc00b;
aud[46828]=16'hc00c;
aud[46829]=16'hc00d;
aud[46830]=16'hc00d;
aud[46831]=16'hc00e;
aud[46832]=16'hc00f;
aud[46833]=16'hc010;
aud[46834]=16'hc011;
aud[46835]=16'hc012;
aud[46836]=16'hc013;
aud[46837]=16'hc014;
aud[46838]=16'hc015;
aud[46839]=16'hc016;
aud[46840]=16'hc018;
aud[46841]=16'hc019;
aud[46842]=16'hc01a;
aud[46843]=16'hc01b;
aud[46844]=16'hc01c;
aud[46845]=16'hc01e;
aud[46846]=16'hc01f;
aud[46847]=16'hc020;
aud[46848]=16'hc022;
aud[46849]=16'hc023;
aud[46850]=16'hc024;
aud[46851]=16'hc026;
aud[46852]=16'hc027;
aud[46853]=16'hc029;
aud[46854]=16'hc02a;
aud[46855]=16'hc02c;
aud[46856]=16'hc02e;
aud[46857]=16'hc02f;
aud[46858]=16'hc031;
aud[46859]=16'hc033;
aud[46860]=16'hc034;
aud[46861]=16'hc036;
aud[46862]=16'hc038;
aud[46863]=16'hc039;
aud[46864]=16'hc03b;
aud[46865]=16'hc03d;
aud[46866]=16'hc03f;
aud[46867]=16'hc041;
aud[46868]=16'hc043;
aud[46869]=16'hc045;
aud[46870]=16'hc047;
aud[46871]=16'hc049;
aud[46872]=16'hc04b;
aud[46873]=16'hc04d;
aud[46874]=16'hc04f;
aud[46875]=16'hc051;
aud[46876]=16'hc053;
aud[46877]=16'hc055;
aud[46878]=16'hc058;
aud[46879]=16'hc05a;
aud[46880]=16'hc05c;
aud[46881]=16'hc05e;
aud[46882]=16'hc061;
aud[46883]=16'hc063;
aud[46884]=16'hc065;
aud[46885]=16'hc068;
aud[46886]=16'hc06a;
aud[46887]=16'hc06d;
aud[46888]=16'hc06f;
aud[46889]=16'hc072;
aud[46890]=16'hc074;
aud[46891]=16'hc077;
aud[46892]=16'hc079;
aud[46893]=16'hc07c;
aud[46894]=16'hc07f;
aud[46895]=16'hc081;
aud[46896]=16'hc084;
aud[46897]=16'hc087;
aud[46898]=16'hc089;
aud[46899]=16'hc08c;
aud[46900]=16'hc08f;
aud[46901]=16'hc092;
aud[46902]=16'hc095;
aud[46903]=16'hc098;
aud[46904]=16'hc09b;
aud[46905]=16'hc09d;
aud[46906]=16'hc0a0;
aud[46907]=16'hc0a3;
aud[46908]=16'hc0a6;
aud[46909]=16'hc0aa;
aud[46910]=16'hc0ad;
aud[46911]=16'hc0b0;
aud[46912]=16'hc0b3;
aud[46913]=16'hc0b6;
aud[46914]=16'hc0b9;
aud[46915]=16'hc0bd;
aud[46916]=16'hc0c0;
aud[46917]=16'hc0c3;
aud[46918]=16'hc0c6;
aud[46919]=16'hc0ca;
aud[46920]=16'hc0cd;
aud[46921]=16'hc0d0;
aud[46922]=16'hc0d4;
aud[46923]=16'hc0d7;
aud[46924]=16'hc0db;
aud[46925]=16'hc0de;
aud[46926]=16'hc0e2;
aud[46927]=16'hc0e5;
aud[46928]=16'hc0e9;
aud[46929]=16'hc0ed;
aud[46930]=16'hc0f0;
aud[46931]=16'hc0f4;
aud[46932]=16'hc0f8;
aud[46933]=16'hc0fb;
aud[46934]=16'hc0ff;
aud[46935]=16'hc103;
aud[46936]=16'hc107;
aud[46937]=16'hc10b;
aud[46938]=16'hc10e;
aud[46939]=16'hc112;
aud[46940]=16'hc116;
aud[46941]=16'hc11a;
aud[46942]=16'hc11e;
aud[46943]=16'hc122;
aud[46944]=16'hc126;
aud[46945]=16'hc12a;
aud[46946]=16'hc12e;
aud[46947]=16'hc133;
aud[46948]=16'hc137;
aud[46949]=16'hc13b;
aud[46950]=16'hc13f;
aud[46951]=16'hc143;
aud[46952]=16'hc147;
aud[46953]=16'hc14c;
aud[46954]=16'hc150;
aud[46955]=16'hc154;
aud[46956]=16'hc159;
aud[46957]=16'hc15d;
aud[46958]=16'hc162;
aud[46959]=16'hc166;
aud[46960]=16'hc16b;
aud[46961]=16'hc16f;
aud[46962]=16'hc174;
aud[46963]=16'hc178;
aud[46964]=16'hc17d;
aud[46965]=16'hc181;
aud[46966]=16'hc186;
aud[46967]=16'hc18b;
aud[46968]=16'hc18f;
aud[46969]=16'hc194;
aud[46970]=16'hc199;
aud[46971]=16'hc19e;
aud[46972]=16'hc1a2;
aud[46973]=16'hc1a7;
aud[46974]=16'hc1ac;
aud[46975]=16'hc1b1;
aud[46976]=16'hc1b6;
aud[46977]=16'hc1bb;
aud[46978]=16'hc1c0;
aud[46979]=16'hc1c5;
aud[46980]=16'hc1ca;
aud[46981]=16'hc1cf;
aud[46982]=16'hc1d4;
aud[46983]=16'hc1d9;
aud[46984]=16'hc1de;
aud[46985]=16'hc1e3;
aud[46986]=16'hc1e8;
aud[46987]=16'hc1ee;
aud[46988]=16'hc1f3;
aud[46989]=16'hc1f8;
aud[46990]=16'hc1fd;
aud[46991]=16'hc203;
aud[46992]=16'hc208;
aud[46993]=16'hc20d;
aud[46994]=16'hc213;
aud[46995]=16'hc218;
aud[46996]=16'hc21e;
aud[46997]=16'hc223;
aud[46998]=16'hc229;
aud[46999]=16'hc22e;
aud[47000]=16'hc234;
aud[47001]=16'hc239;
aud[47002]=16'hc23f;
aud[47003]=16'hc245;
aud[47004]=16'hc24a;
aud[47005]=16'hc250;
aud[47006]=16'hc256;
aud[47007]=16'hc25c;
aud[47008]=16'hc261;
aud[47009]=16'hc267;
aud[47010]=16'hc26d;
aud[47011]=16'hc273;
aud[47012]=16'hc279;
aud[47013]=16'hc27f;
aud[47014]=16'hc285;
aud[47015]=16'hc28b;
aud[47016]=16'hc291;
aud[47017]=16'hc297;
aud[47018]=16'hc29d;
aud[47019]=16'hc2a3;
aud[47020]=16'hc2a9;
aud[47021]=16'hc2af;
aud[47022]=16'hc2b5;
aud[47023]=16'hc2bb;
aud[47024]=16'hc2c1;
aud[47025]=16'hc2c8;
aud[47026]=16'hc2ce;
aud[47027]=16'hc2d4;
aud[47028]=16'hc2db;
aud[47029]=16'hc2e1;
aud[47030]=16'hc2e7;
aud[47031]=16'hc2ee;
aud[47032]=16'hc2f4;
aud[47033]=16'hc2fb;
aud[47034]=16'hc301;
aud[47035]=16'hc308;
aud[47036]=16'hc30e;
aud[47037]=16'hc315;
aud[47038]=16'hc31b;
aud[47039]=16'hc322;
aud[47040]=16'hc329;
aud[47041]=16'hc32f;
aud[47042]=16'hc336;
aud[47043]=16'hc33d;
aud[47044]=16'hc343;
aud[47045]=16'hc34a;
aud[47046]=16'hc351;
aud[47047]=16'hc358;
aud[47048]=16'hc35f;
aud[47049]=16'hc365;
aud[47050]=16'hc36c;
aud[47051]=16'hc373;
aud[47052]=16'hc37a;
aud[47053]=16'hc381;
aud[47054]=16'hc388;
aud[47055]=16'hc38f;
aud[47056]=16'hc396;
aud[47057]=16'hc39d;
aud[47058]=16'hc3a5;
aud[47059]=16'hc3ac;
aud[47060]=16'hc3b3;
aud[47061]=16'hc3ba;
aud[47062]=16'hc3c1;
aud[47063]=16'hc3c9;
aud[47064]=16'hc3d0;
aud[47065]=16'hc3d7;
aud[47066]=16'hc3df;
aud[47067]=16'hc3e6;
aud[47068]=16'hc3ed;
aud[47069]=16'hc3f5;
aud[47070]=16'hc3fc;
aud[47071]=16'hc404;
aud[47072]=16'hc40b;
aud[47073]=16'hc413;
aud[47074]=16'hc41a;
aud[47075]=16'hc422;
aud[47076]=16'hc429;
aud[47077]=16'hc431;
aud[47078]=16'hc439;
aud[47079]=16'hc440;
aud[47080]=16'hc448;
aud[47081]=16'hc450;
aud[47082]=16'hc457;
aud[47083]=16'hc45f;
aud[47084]=16'hc467;
aud[47085]=16'hc46f;
aud[47086]=16'hc477;
aud[47087]=16'hc47f;
aud[47088]=16'hc486;
aud[47089]=16'hc48e;
aud[47090]=16'hc496;
aud[47091]=16'hc49e;
aud[47092]=16'hc4a6;
aud[47093]=16'hc4ae;
aud[47094]=16'hc4b6;
aud[47095]=16'hc4bf;
aud[47096]=16'hc4c7;
aud[47097]=16'hc4cf;
aud[47098]=16'hc4d7;
aud[47099]=16'hc4df;
aud[47100]=16'hc4e7;
aud[47101]=16'hc4f0;
aud[47102]=16'hc4f8;
aud[47103]=16'hc500;
aud[47104]=16'hc509;
aud[47105]=16'hc511;
aud[47106]=16'hc519;
aud[47107]=16'hc522;
aud[47108]=16'hc52a;
aud[47109]=16'hc533;
aud[47110]=16'hc53b;
aud[47111]=16'hc544;
aud[47112]=16'hc54c;
aud[47113]=16'hc555;
aud[47114]=16'hc55d;
aud[47115]=16'hc566;
aud[47116]=16'hc56e;
aud[47117]=16'hc577;
aud[47118]=16'hc580;
aud[47119]=16'hc588;
aud[47120]=16'hc591;
aud[47121]=16'hc59a;
aud[47122]=16'hc5a3;
aud[47123]=16'hc5ac;
aud[47124]=16'hc5b4;
aud[47125]=16'hc5bd;
aud[47126]=16'hc5c6;
aud[47127]=16'hc5cf;
aud[47128]=16'hc5d8;
aud[47129]=16'hc5e1;
aud[47130]=16'hc5ea;
aud[47131]=16'hc5f3;
aud[47132]=16'hc5fc;
aud[47133]=16'hc605;
aud[47134]=16'hc60e;
aud[47135]=16'hc617;
aud[47136]=16'hc620;
aud[47137]=16'hc62a;
aud[47138]=16'hc633;
aud[47139]=16'hc63c;
aud[47140]=16'hc645;
aud[47141]=16'hc64f;
aud[47142]=16'hc658;
aud[47143]=16'hc661;
aud[47144]=16'hc66b;
aud[47145]=16'hc674;
aud[47146]=16'hc67d;
aud[47147]=16'hc687;
aud[47148]=16'hc690;
aud[47149]=16'hc69a;
aud[47150]=16'hc6a3;
aud[47151]=16'hc6ad;
aud[47152]=16'hc6b6;
aud[47153]=16'hc6c0;
aud[47154]=16'hc6c9;
aud[47155]=16'hc6d3;
aud[47156]=16'hc6dd;
aud[47157]=16'hc6e6;
aud[47158]=16'hc6f0;
aud[47159]=16'hc6fa;
aud[47160]=16'hc703;
aud[47161]=16'hc70d;
aud[47162]=16'hc717;
aud[47163]=16'hc721;
aud[47164]=16'hc72b;
aud[47165]=16'hc735;
aud[47166]=16'hc73f;
aud[47167]=16'hc748;
aud[47168]=16'hc752;
aud[47169]=16'hc75c;
aud[47170]=16'hc766;
aud[47171]=16'hc770;
aud[47172]=16'hc77a;
aud[47173]=16'hc785;
aud[47174]=16'hc78f;
aud[47175]=16'hc799;
aud[47176]=16'hc7a3;
aud[47177]=16'hc7ad;
aud[47178]=16'hc7b7;
aud[47179]=16'hc7c1;
aud[47180]=16'hc7cc;
aud[47181]=16'hc7d6;
aud[47182]=16'hc7e0;
aud[47183]=16'hc7eb;
aud[47184]=16'hc7f5;
aud[47185]=16'hc7ff;
aud[47186]=16'hc80a;
aud[47187]=16'hc814;
aud[47188]=16'hc81f;
aud[47189]=16'hc829;
aud[47190]=16'hc834;
aud[47191]=16'hc83e;
aud[47192]=16'hc849;
aud[47193]=16'hc853;
aud[47194]=16'hc85e;
aud[47195]=16'hc868;
aud[47196]=16'hc873;
aud[47197]=16'hc87e;
aud[47198]=16'hc888;
aud[47199]=16'hc893;
aud[47200]=16'hc89e;
aud[47201]=16'hc8a9;
aud[47202]=16'hc8b3;
aud[47203]=16'hc8be;
aud[47204]=16'hc8c9;
aud[47205]=16'hc8d4;
aud[47206]=16'hc8df;
aud[47207]=16'hc8ea;
aud[47208]=16'hc8f5;
aud[47209]=16'hc8ff;
aud[47210]=16'hc90a;
aud[47211]=16'hc915;
aud[47212]=16'hc920;
aud[47213]=16'hc92c;
aud[47214]=16'hc937;
aud[47215]=16'hc942;
aud[47216]=16'hc94d;
aud[47217]=16'hc958;
aud[47218]=16'hc963;
aud[47219]=16'hc96e;
aud[47220]=16'hc97a;
aud[47221]=16'hc985;
aud[47222]=16'hc990;
aud[47223]=16'hc99b;
aud[47224]=16'hc9a7;
aud[47225]=16'hc9b2;
aud[47226]=16'hc9bd;
aud[47227]=16'hc9c9;
aud[47228]=16'hc9d4;
aud[47229]=16'hc9e0;
aud[47230]=16'hc9eb;
aud[47231]=16'hc9f7;
aud[47232]=16'hca02;
aud[47233]=16'hca0e;
aud[47234]=16'hca19;
aud[47235]=16'hca25;
aud[47236]=16'hca30;
aud[47237]=16'hca3c;
aud[47238]=16'hca48;
aud[47239]=16'hca53;
aud[47240]=16'hca5f;
aud[47241]=16'hca6b;
aud[47242]=16'hca76;
aud[47243]=16'hca82;
aud[47244]=16'hca8e;
aud[47245]=16'hca9a;
aud[47246]=16'hcaa6;
aud[47247]=16'hcab1;
aud[47248]=16'hcabd;
aud[47249]=16'hcac9;
aud[47250]=16'hcad5;
aud[47251]=16'hcae1;
aud[47252]=16'hcaed;
aud[47253]=16'hcaf9;
aud[47254]=16'hcb05;
aud[47255]=16'hcb11;
aud[47256]=16'hcb1d;
aud[47257]=16'hcb29;
aud[47258]=16'hcb35;
aud[47259]=16'hcb42;
aud[47260]=16'hcb4e;
aud[47261]=16'hcb5a;
aud[47262]=16'hcb66;
aud[47263]=16'hcb72;
aud[47264]=16'hcb7f;
aud[47265]=16'hcb8b;
aud[47266]=16'hcb97;
aud[47267]=16'hcba3;
aud[47268]=16'hcbb0;
aud[47269]=16'hcbbc;
aud[47270]=16'hcbc9;
aud[47271]=16'hcbd5;
aud[47272]=16'hcbe1;
aud[47273]=16'hcbee;
aud[47274]=16'hcbfa;
aud[47275]=16'hcc07;
aud[47276]=16'hcc13;
aud[47277]=16'hcc20;
aud[47278]=16'hcc2c;
aud[47279]=16'hcc39;
aud[47280]=16'hcc46;
aud[47281]=16'hcc52;
aud[47282]=16'hcc5f;
aud[47283]=16'hcc6c;
aud[47284]=16'hcc78;
aud[47285]=16'hcc85;
aud[47286]=16'hcc92;
aud[47287]=16'hcc9f;
aud[47288]=16'hccab;
aud[47289]=16'hccb8;
aud[47290]=16'hccc5;
aud[47291]=16'hccd2;
aud[47292]=16'hccdf;
aud[47293]=16'hccec;
aud[47294]=16'hccf9;
aud[47295]=16'hcd06;
aud[47296]=16'hcd13;
aud[47297]=16'hcd20;
aud[47298]=16'hcd2d;
aud[47299]=16'hcd3a;
aud[47300]=16'hcd47;
aud[47301]=16'hcd54;
aud[47302]=16'hcd61;
aud[47303]=16'hcd6e;
aud[47304]=16'hcd7b;
aud[47305]=16'hcd88;
aud[47306]=16'hcd96;
aud[47307]=16'hcda3;
aud[47308]=16'hcdb0;
aud[47309]=16'hcdbd;
aud[47310]=16'hcdcb;
aud[47311]=16'hcdd8;
aud[47312]=16'hcde5;
aud[47313]=16'hcdf3;
aud[47314]=16'hce00;
aud[47315]=16'hce0d;
aud[47316]=16'hce1b;
aud[47317]=16'hce28;
aud[47318]=16'hce36;
aud[47319]=16'hce43;
aud[47320]=16'hce51;
aud[47321]=16'hce5e;
aud[47322]=16'hce6c;
aud[47323]=16'hce79;
aud[47324]=16'hce87;
aud[47325]=16'hce95;
aud[47326]=16'hcea2;
aud[47327]=16'hceb0;
aud[47328]=16'hcebe;
aud[47329]=16'hcecb;
aud[47330]=16'hced9;
aud[47331]=16'hcee7;
aud[47332]=16'hcef5;
aud[47333]=16'hcf02;
aud[47334]=16'hcf10;
aud[47335]=16'hcf1e;
aud[47336]=16'hcf2c;
aud[47337]=16'hcf3a;
aud[47338]=16'hcf48;
aud[47339]=16'hcf56;
aud[47340]=16'hcf63;
aud[47341]=16'hcf71;
aud[47342]=16'hcf7f;
aud[47343]=16'hcf8d;
aud[47344]=16'hcf9b;
aud[47345]=16'hcfa9;
aud[47346]=16'hcfb8;
aud[47347]=16'hcfc6;
aud[47348]=16'hcfd4;
aud[47349]=16'hcfe2;
aud[47350]=16'hcff0;
aud[47351]=16'hcffe;
aud[47352]=16'hd00c;
aud[47353]=16'hd01b;
aud[47354]=16'hd029;
aud[47355]=16'hd037;
aud[47356]=16'hd045;
aud[47357]=16'hd054;
aud[47358]=16'hd062;
aud[47359]=16'hd070;
aud[47360]=16'hd07f;
aud[47361]=16'hd08d;
aud[47362]=16'hd09b;
aud[47363]=16'hd0aa;
aud[47364]=16'hd0b8;
aud[47365]=16'hd0c7;
aud[47366]=16'hd0d5;
aud[47367]=16'hd0e4;
aud[47368]=16'hd0f2;
aud[47369]=16'hd101;
aud[47370]=16'hd10f;
aud[47371]=16'hd11e;
aud[47372]=16'hd12d;
aud[47373]=16'hd13b;
aud[47374]=16'hd14a;
aud[47375]=16'hd159;
aud[47376]=16'hd167;
aud[47377]=16'hd176;
aud[47378]=16'hd185;
aud[47379]=16'hd193;
aud[47380]=16'hd1a2;
aud[47381]=16'hd1b1;
aud[47382]=16'hd1c0;
aud[47383]=16'hd1cf;
aud[47384]=16'hd1de;
aud[47385]=16'hd1ec;
aud[47386]=16'hd1fb;
aud[47387]=16'hd20a;
aud[47388]=16'hd219;
aud[47389]=16'hd228;
aud[47390]=16'hd237;
aud[47391]=16'hd246;
aud[47392]=16'hd255;
aud[47393]=16'hd264;
aud[47394]=16'hd273;
aud[47395]=16'hd282;
aud[47396]=16'hd291;
aud[47397]=16'hd2a0;
aud[47398]=16'hd2b0;
aud[47399]=16'hd2bf;
aud[47400]=16'hd2ce;
aud[47401]=16'hd2dd;
aud[47402]=16'hd2ec;
aud[47403]=16'hd2fc;
aud[47404]=16'hd30b;
aud[47405]=16'hd31a;
aud[47406]=16'hd329;
aud[47407]=16'hd339;
aud[47408]=16'hd348;
aud[47409]=16'hd357;
aud[47410]=16'hd367;
aud[47411]=16'hd376;
aud[47412]=16'hd386;
aud[47413]=16'hd395;
aud[47414]=16'hd3a4;
aud[47415]=16'hd3b4;
aud[47416]=16'hd3c3;
aud[47417]=16'hd3d3;
aud[47418]=16'hd3e2;
aud[47419]=16'hd3f2;
aud[47420]=16'hd402;
aud[47421]=16'hd411;
aud[47422]=16'hd421;
aud[47423]=16'hd430;
aud[47424]=16'hd440;
aud[47425]=16'hd450;
aud[47426]=16'hd45f;
aud[47427]=16'hd46f;
aud[47428]=16'hd47f;
aud[47429]=16'hd48f;
aud[47430]=16'hd49e;
aud[47431]=16'hd4ae;
aud[47432]=16'hd4be;
aud[47433]=16'hd4ce;
aud[47434]=16'hd4de;
aud[47435]=16'hd4ed;
aud[47436]=16'hd4fd;
aud[47437]=16'hd50d;
aud[47438]=16'hd51d;
aud[47439]=16'hd52d;
aud[47440]=16'hd53d;
aud[47441]=16'hd54d;
aud[47442]=16'hd55d;
aud[47443]=16'hd56d;
aud[47444]=16'hd57d;
aud[47445]=16'hd58d;
aud[47446]=16'hd59d;
aud[47447]=16'hd5ad;
aud[47448]=16'hd5bd;
aud[47449]=16'hd5cd;
aud[47450]=16'hd5dd;
aud[47451]=16'hd5ee;
aud[47452]=16'hd5fe;
aud[47453]=16'hd60e;
aud[47454]=16'hd61e;
aud[47455]=16'hd62e;
aud[47456]=16'hd63f;
aud[47457]=16'hd64f;
aud[47458]=16'hd65f;
aud[47459]=16'hd66f;
aud[47460]=16'hd680;
aud[47461]=16'hd690;
aud[47462]=16'hd6a0;
aud[47463]=16'hd6b1;
aud[47464]=16'hd6c1;
aud[47465]=16'hd6d2;
aud[47466]=16'hd6e2;
aud[47467]=16'hd6f2;
aud[47468]=16'hd703;
aud[47469]=16'hd713;
aud[47470]=16'hd724;
aud[47471]=16'hd734;
aud[47472]=16'hd745;
aud[47473]=16'hd756;
aud[47474]=16'hd766;
aud[47475]=16'hd777;
aud[47476]=16'hd787;
aud[47477]=16'hd798;
aud[47478]=16'hd7a9;
aud[47479]=16'hd7b9;
aud[47480]=16'hd7ca;
aud[47481]=16'hd7db;
aud[47482]=16'hd7eb;
aud[47483]=16'hd7fc;
aud[47484]=16'hd80d;
aud[47485]=16'hd81e;
aud[47486]=16'hd82e;
aud[47487]=16'hd83f;
aud[47488]=16'hd850;
aud[47489]=16'hd861;
aud[47490]=16'hd872;
aud[47491]=16'hd882;
aud[47492]=16'hd893;
aud[47493]=16'hd8a4;
aud[47494]=16'hd8b5;
aud[47495]=16'hd8c6;
aud[47496]=16'hd8d7;
aud[47497]=16'hd8e8;
aud[47498]=16'hd8f9;
aud[47499]=16'hd90a;
aud[47500]=16'hd91b;
aud[47501]=16'hd92c;
aud[47502]=16'hd93d;
aud[47503]=16'hd94e;
aud[47504]=16'hd95f;
aud[47505]=16'hd970;
aud[47506]=16'hd982;
aud[47507]=16'hd993;
aud[47508]=16'hd9a4;
aud[47509]=16'hd9b5;
aud[47510]=16'hd9c6;
aud[47511]=16'hd9d7;
aud[47512]=16'hd9e9;
aud[47513]=16'hd9fa;
aud[47514]=16'hda0b;
aud[47515]=16'hda1c;
aud[47516]=16'hda2e;
aud[47517]=16'hda3f;
aud[47518]=16'hda50;
aud[47519]=16'hda62;
aud[47520]=16'hda73;
aud[47521]=16'hda84;
aud[47522]=16'hda96;
aud[47523]=16'hdaa7;
aud[47524]=16'hdab9;
aud[47525]=16'hdaca;
aud[47526]=16'hdadc;
aud[47527]=16'hdaed;
aud[47528]=16'hdaff;
aud[47529]=16'hdb10;
aud[47530]=16'hdb22;
aud[47531]=16'hdb33;
aud[47532]=16'hdb45;
aud[47533]=16'hdb56;
aud[47534]=16'hdb68;
aud[47535]=16'hdb79;
aud[47536]=16'hdb8b;
aud[47537]=16'hdb9d;
aud[47538]=16'hdbae;
aud[47539]=16'hdbc0;
aud[47540]=16'hdbd2;
aud[47541]=16'hdbe3;
aud[47542]=16'hdbf5;
aud[47543]=16'hdc07;
aud[47544]=16'hdc19;
aud[47545]=16'hdc2a;
aud[47546]=16'hdc3c;
aud[47547]=16'hdc4e;
aud[47548]=16'hdc60;
aud[47549]=16'hdc72;
aud[47550]=16'hdc83;
aud[47551]=16'hdc95;
aud[47552]=16'hdca7;
aud[47553]=16'hdcb9;
aud[47554]=16'hdccb;
aud[47555]=16'hdcdd;
aud[47556]=16'hdcef;
aud[47557]=16'hdd01;
aud[47558]=16'hdd13;
aud[47559]=16'hdd25;
aud[47560]=16'hdd37;
aud[47561]=16'hdd49;
aud[47562]=16'hdd5b;
aud[47563]=16'hdd6d;
aud[47564]=16'hdd7f;
aud[47565]=16'hdd91;
aud[47566]=16'hdda3;
aud[47567]=16'hddb5;
aud[47568]=16'hddc7;
aud[47569]=16'hddd9;
aud[47570]=16'hddeb;
aud[47571]=16'hddfe;
aud[47572]=16'hde10;
aud[47573]=16'hde22;
aud[47574]=16'hde34;
aud[47575]=16'hde46;
aud[47576]=16'hde59;
aud[47577]=16'hde6b;
aud[47578]=16'hde7d;
aud[47579]=16'hde8f;
aud[47580]=16'hdea2;
aud[47581]=16'hdeb4;
aud[47582]=16'hdec6;
aud[47583]=16'hded9;
aud[47584]=16'hdeeb;
aud[47585]=16'hdefd;
aud[47586]=16'hdf10;
aud[47587]=16'hdf22;
aud[47588]=16'hdf35;
aud[47589]=16'hdf47;
aud[47590]=16'hdf59;
aud[47591]=16'hdf6c;
aud[47592]=16'hdf7e;
aud[47593]=16'hdf91;
aud[47594]=16'hdfa3;
aud[47595]=16'hdfb6;
aud[47596]=16'hdfc8;
aud[47597]=16'hdfdb;
aud[47598]=16'hdfed;
aud[47599]=16'he000;
aud[47600]=16'he013;
aud[47601]=16'he025;
aud[47602]=16'he038;
aud[47603]=16'he04a;
aud[47604]=16'he05d;
aud[47605]=16'he070;
aud[47606]=16'he082;
aud[47607]=16'he095;
aud[47608]=16'he0a8;
aud[47609]=16'he0ba;
aud[47610]=16'he0cd;
aud[47611]=16'he0e0;
aud[47612]=16'he0f3;
aud[47613]=16'he105;
aud[47614]=16'he118;
aud[47615]=16'he12b;
aud[47616]=16'he13e;
aud[47617]=16'he151;
aud[47618]=16'he163;
aud[47619]=16'he176;
aud[47620]=16'he189;
aud[47621]=16'he19c;
aud[47622]=16'he1af;
aud[47623]=16'he1c2;
aud[47624]=16'he1d5;
aud[47625]=16'he1e8;
aud[47626]=16'he1fa;
aud[47627]=16'he20d;
aud[47628]=16'he220;
aud[47629]=16'he233;
aud[47630]=16'he246;
aud[47631]=16'he259;
aud[47632]=16'he26c;
aud[47633]=16'he27f;
aud[47634]=16'he292;
aud[47635]=16'he2a5;
aud[47636]=16'he2b9;
aud[47637]=16'he2cc;
aud[47638]=16'he2df;
aud[47639]=16'he2f2;
aud[47640]=16'he305;
aud[47641]=16'he318;
aud[47642]=16'he32b;
aud[47643]=16'he33e;
aud[47644]=16'he352;
aud[47645]=16'he365;
aud[47646]=16'he378;
aud[47647]=16'he38b;
aud[47648]=16'he39e;
aud[47649]=16'he3b2;
aud[47650]=16'he3c5;
aud[47651]=16'he3d8;
aud[47652]=16'he3eb;
aud[47653]=16'he3ff;
aud[47654]=16'he412;
aud[47655]=16'he425;
aud[47656]=16'he438;
aud[47657]=16'he44c;
aud[47658]=16'he45f;
aud[47659]=16'he473;
aud[47660]=16'he486;
aud[47661]=16'he499;
aud[47662]=16'he4ad;
aud[47663]=16'he4c0;
aud[47664]=16'he4d3;
aud[47665]=16'he4e7;
aud[47666]=16'he4fa;
aud[47667]=16'he50e;
aud[47668]=16'he521;
aud[47669]=16'he535;
aud[47670]=16'he548;
aud[47671]=16'he55c;
aud[47672]=16'he56f;
aud[47673]=16'he583;
aud[47674]=16'he596;
aud[47675]=16'he5aa;
aud[47676]=16'he5bd;
aud[47677]=16'he5d1;
aud[47678]=16'he5e4;
aud[47679]=16'he5f8;
aud[47680]=16'he60c;
aud[47681]=16'he61f;
aud[47682]=16'he633;
aud[47683]=16'he646;
aud[47684]=16'he65a;
aud[47685]=16'he66e;
aud[47686]=16'he681;
aud[47687]=16'he695;
aud[47688]=16'he6a9;
aud[47689]=16'he6bd;
aud[47690]=16'he6d0;
aud[47691]=16'he6e4;
aud[47692]=16'he6f8;
aud[47693]=16'he70b;
aud[47694]=16'he71f;
aud[47695]=16'he733;
aud[47696]=16'he747;
aud[47697]=16'he75b;
aud[47698]=16'he76e;
aud[47699]=16'he782;
aud[47700]=16'he796;
aud[47701]=16'he7aa;
aud[47702]=16'he7be;
aud[47703]=16'he7d1;
aud[47704]=16'he7e5;
aud[47705]=16'he7f9;
aud[47706]=16'he80d;
aud[47707]=16'he821;
aud[47708]=16'he835;
aud[47709]=16'he849;
aud[47710]=16'he85d;
aud[47711]=16'he871;
aud[47712]=16'he885;
aud[47713]=16'he899;
aud[47714]=16'he8ad;
aud[47715]=16'he8c0;
aud[47716]=16'he8d4;
aud[47717]=16'he8e8;
aud[47718]=16'he8fc;
aud[47719]=16'he910;
aud[47720]=16'he925;
aud[47721]=16'he939;
aud[47722]=16'he94d;
aud[47723]=16'he961;
aud[47724]=16'he975;
aud[47725]=16'he989;
aud[47726]=16'he99d;
aud[47727]=16'he9b1;
aud[47728]=16'he9c5;
aud[47729]=16'he9d9;
aud[47730]=16'he9ed;
aud[47731]=16'hea01;
aud[47732]=16'hea16;
aud[47733]=16'hea2a;
aud[47734]=16'hea3e;
aud[47735]=16'hea52;
aud[47736]=16'hea66;
aud[47737]=16'hea7a;
aud[47738]=16'hea8f;
aud[47739]=16'heaa3;
aud[47740]=16'heab7;
aud[47741]=16'heacb;
aud[47742]=16'heae0;
aud[47743]=16'heaf4;
aud[47744]=16'heb08;
aud[47745]=16'heb1c;
aud[47746]=16'heb31;
aud[47747]=16'heb45;
aud[47748]=16'heb59;
aud[47749]=16'heb6e;
aud[47750]=16'heb82;
aud[47751]=16'heb96;
aud[47752]=16'hebab;
aud[47753]=16'hebbf;
aud[47754]=16'hebd3;
aud[47755]=16'hebe8;
aud[47756]=16'hebfc;
aud[47757]=16'hec10;
aud[47758]=16'hec25;
aud[47759]=16'hec39;
aud[47760]=16'hec4d;
aud[47761]=16'hec62;
aud[47762]=16'hec76;
aud[47763]=16'hec8b;
aud[47764]=16'hec9f;
aud[47765]=16'hecb4;
aud[47766]=16'hecc8;
aud[47767]=16'hecdd;
aud[47768]=16'hecf1;
aud[47769]=16'hed05;
aud[47770]=16'hed1a;
aud[47771]=16'hed2e;
aud[47772]=16'hed43;
aud[47773]=16'hed57;
aud[47774]=16'hed6c;
aud[47775]=16'hed81;
aud[47776]=16'hed95;
aud[47777]=16'hedaa;
aud[47778]=16'hedbe;
aud[47779]=16'hedd3;
aud[47780]=16'hede7;
aud[47781]=16'hedfc;
aud[47782]=16'hee10;
aud[47783]=16'hee25;
aud[47784]=16'hee3a;
aud[47785]=16'hee4e;
aud[47786]=16'hee63;
aud[47787]=16'hee77;
aud[47788]=16'hee8c;
aud[47789]=16'heea1;
aud[47790]=16'heeb5;
aud[47791]=16'heeca;
aud[47792]=16'heedf;
aud[47793]=16'heef3;
aud[47794]=16'hef08;
aud[47795]=16'hef1d;
aud[47796]=16'hef31;
aud[47797]=16'hef46;
aud[47798]=16'hef5b;
aud[47799]=16'hef70;
aud[47800]=16'hef84;
aud[47801]=16'hef99;
aud[47802]=16'hefae;
aud[47803]=16'hefc2;
aud[47804]=16'hefd7;
aud[47805]=16'hefec;
aud[47806]=16'hf001;
aud[47807]=16'hf015;
aud[47808]=16'hf02a;
aud[47809]=16'hf03f;
aud[47810]=16'hf054;
aud[47811]=16'hf069;
aud[47812]=16'hf07d;
aud[47813]=16'hf092;
aud[47814]=16'hf0a7;
aud[47815]=16'hf0bc;
aud[47816]=16'hf0d1;
aud[47817]=16'hf0e6;
aud[47818]=16'hf0fa;
aud[47819]=16'hf10f;
aud[47820]=16'hf124;
aud[47821]=16'hf139;
aud[47822]=16'hf14e;
aud[47823]=16'hf163;
aud[47824]=16'hf178;
aud[47825]=16'hf18c;
aud[47826]=16'hf1a1;
aud[47827]=16'hf1b6;
aud[47828]=16'hf1cb;
aud[47829]=16'hf1e0;
aud[47830]=16'hf1f5;
aud[47831]=16'hf20a;
aud[47832]=16'hf21f;
aud[47833]=16'hf234;
aud[47834]=16'hf249;
aud[47835]=16'hf25e;
aud[47836]=16'hf273;
aud[47837]=16'hf288;
aud[47838]=16'hf29d;
aud[47839]=16'hf2b2;
aud[47840]=16'hf2c7;
aud[47841]=16'hf2dc;
aud[47842]=16'hf2f1;
aud[47843]=16'hf306;
aud[47844]=16'hf31b;
aud[47845]=16'hf330;
aud[47846]=16'hf345;
aud[47847]=16'hf35a;
aud[47848]=16'hf36f;
aud[47849]=16'hf384;
aud[47850]=16'hf399;
aud[47851]=16'hf3ae;
aud[47852]=16'hf3c3;
aud[47853]=16'hf3d8;
aud[47854]=16'hf3ed;
aud[47855]=16'hf402;
aud[47856]=16'hf417;
aud[47857]=16'hf42c;
aud[47858]=16'hf441;
aud[47859]=16'hf456;
aud[47860]=16'hf46b;
aud[47861]=16'hf480;
aud[47862]=16'hf496;
aud[47863]=16'hf4ab;
aud[47864]=16'hf4c0;
aud[47865]=16'hf4d5;
aud[47866]=16'hf4ea;
aud[47867]=16'hf4ff;
aud[47868]=16'hf514;
aud[47869]=16'hf529;
aud[47870]=16'hf53f;
aud[47871]=16'hf554;
aud[47872]=16'hf569;
aud[47873]=16'hf57e;
aud[47874]=16'hf593;
aud[47875]=16'hf5a8;
aud[47876]=16'hf5bd;
aud[47877]=16'hf5d3;
aud[47878]=16'hf5e8;
aud[47879]=16'hf5fd;
aud[47880]=16'hf612;
aud[47881]=16'hf627;
aud[47882]=16'hf63d;
aud[47883]=16'hf652;
aud[47884]=16'hf667;
aud[47885]=16'hf67c;
aud[47886]=16'hf691;
aud[47887]=16'hf6a7;
aud[47888]=16'hf6bc;
aud[47889]=16'hf6d1;
aud[47890]=16'hf6e6;
aud[47891]=16'hf6fb;
aud[47892]=16'hf711;
aud[47893]=16'hf726;
aud[47894]=16'hf73b;
aud[47895]=16'hf750;
aud[47896]=16'hf766;
aud[47897]=16'hf77b;
aud[47898]=16'hf790;
aud[47899]=16'hf7a5;
aud[47900]=16'hf7bb;
aud[47901]=16'hf7d0;
aud[47902]=16'hf7e5;
aud[47903]=16'hf7fb;
aud[47904]=16'hf810;
aud[47905]=16'hf825;
aud[47906]=16'hf83a;
aud[47907]=16'hf850;
aud[47908]=16'hf865;
aud[47909]=16'hf87a;
aud[47910]=16'hf890;
aud[47911]=16'hf8a5;
aud[47912]=16'hf8ba;
aud[47913]=16'hf8cf;
aud[47914]=16'hf8e5;
aud[47915]=16'hf8fa;
aud[47916]=16'hf90f;
aud[47917]=16'hf925;
aud[47918]=16'hf93a;
aud[47919]=16'hf94f;
aud[47920]=16'hf965;
aud[47921]=16'hf97a;
aud[47922]=16'hf98f;
aud[47923]=16'hf9a5;
aud[47924]=16'hf9ba;
aud[47925]=16'hf9cf;
aud[47926]=16'hf9e5;
aud[47927]=16'hf9fa;
aud[47928]=16'hfa0f;
aud[47929]=16'hfa25;
aud[47930]=16'hfa3a;
aud[47931]=16'hfa50;
aud[47932]=16'hfa65;
aud[47933]=16'hfa7a;
aud[47934]=16'hfa90;
aud[47935]=16'hfaa5;
aud[47936]=16'hfaba;
aud[47937]=16'hfad0;
aud[47938]=16'hfae5;
aud[47939]=16'hfafb;
aud[47940]=16'hfb10;
aud[47941]=16'hfb25;
aud[47942]=16'hfb3b;
aud[47943]=16'hfb50;
aud[47944]=16'hfb65;
aud[47945]=16'hfb7b;
aud[47946]=16'hfb90;
aud[47947]=16'hfba6;
aud[47948]=16'hfbbb;
aud[47949]=16'hfbd0;
aud[47950]=16'hfbe6;
aud[47951]=16'hfbfb;
aud[47952]=16'hfc11;
aud[47953]=16'hfc26;
aud[47954]=16'hfc3b;
aud[47955]=16'hfc51;
aud[47956]=16'hfc66;
aud[47957]=16'hfc7c;
aud[47958]=16'hfc91;
aud[47959]=16'hfca7;
aud[47960]=16'hfcbc;
aud[47961]=16'hfcd1;
aud[47962]=16'hfce7;
aud[47963]=16'hfcfc;
aud[47964]=16'hfd12;
aud[47965]=16'hfd27;
aud[47966]=16'hfd3c;
aud[47967]=16'hfd52;
aud[47968]=16'hfd67;
aud[47969]=16'hfd7d;
aud[47970]=16'hfd92;
aud[47971]=16'hfda8;
aud[47972]=16'hfdbd;
aud[47973]=16'hfdd2;
aud[47974]=16'hfde8;
aud[47975]=16'hfdfd;
aud[47976]=16'hfe13;
aud[47977]=16'hfe28;
aud[47978]=16'hfe3e;
aud[47979]=16'hfe53;
aud[47980]=16'hfe69;
aud[47981]=16'hfe7e;
aud[47982]=16'hfe93;
aud[47983]=16'hfea9;
aud[47984]=16'hfebe;
aud[47985]=16'hfed4;
aud[47986]=16'hfee9;
aud[47987]=16'hfeff;
aud[47988]=16'hff14;
aud[47989]=16'hff2a;
aud[47990]=16'hff3f;
aud[47991]=16'hff54;
aud[47992]=16'hff6a;
aud[47993]=16'hff7f;
aud[47994]=16'hff95;
aud[47995]=16'hffaa;
aud[47996]=16'hffc0;
aud[47997]=16'hffd5;
aud[47998]=16'hffeb;
aud[47999]=16'h0;
aud[48000]=16'h15;
aud[48001]=16'h2b;
aud[48002]=16'h40;
aud[48003]=16'h56;
aud[48004]=16'h6b;
aud[48005]=16'h81;
aud[48006]=16'h96;
aud[48007]=16'hac;
aud[48008]=16'hc1;
aud[48009]=16'hd6;
aud[48010]=16'hec;
aud[48011]=16'h101;
aud[48012]=16'h117;
aud[48013]=16'h12c;
aud[48014]=16'h142;
aud[48015]=16'h157;
aud[48016]=16'h16d;
aud[48017]=16'h182;
aud[48018]=16'h197;
aud[48019]=16'h1ad;
aud[48020]=16'h1c2;
aud[48021]=16'h1d8;
aud[48022]=16'h1ed;
aud[48023]=16'h203;
aud[48024]=16'h218;
aud[48025]=16'h22e;
aud[48026]=16'h243;
aud[48027]=16'h258;
aud[48028]=16'h26e;
aud[48029]=16'h283;
aud[48030]=16'h299;
aud[48031]=16'h2ae;
aud[48032]=16'h2c4;
aud[48033]=16'h2d9;
aud[48034]=16'h2ee;
aud[48035]=16'h304;
aud[48036]=16'h319;
aud[48037]=16'h32f;
aud[48038]=16'h344;
aud[48039]=16'h359;
aud[48040]=16'h36f;
aud[48041]=16'h384;
aud[48042]=16'h39a;
aud[48043]=16'h3af;
aud[48044]=16'h3c5;
aud[48045]=16'h3da;
aud[48046]=16'h3ef;
aud[48047]=16'h405;
aud[48048]=16'h41a;
aud[48049]=16'h430;
aud[48050]=16'h445;
aud[48051]=16'h45a;
aud[48052]=16'h470;
aud[48053]=16'h485;
aud[48054]=16'h49b;
aud[48055]=16'h4b0;
aud[48056]=16'h4c5;
aud[48057]=16'h4db;
aud[48058]=16'h4f0;
aud[48059]=16'h505;
aud[48060]=16'h51b;
aud[48061]=16'h530;
aud[48062]=16'h546;
aud[48063]=16'h55b;
aud[48064]=16'h570;
aud[48065]=16'h586;
aud[48066]=16'h59b;
aud[48067]=16'h5b0;
aud[48068]=16'h5c6;
aud[48069]=16'h5db;
aud[48070]=16'h5f1;
aud[48071]=16'h606;
aud[48072]=16'h61b;
aud[48073]=16'h631;
aud[48074]=16'h646;
aud[48075]=16'h65b;
aud[48076]=16'h671;
aud[48077]=16'h686;
aud[48078]=16'h69b;
aud[48079]=16'h6b1;
aud[48080]=16'h6c6;
aud[48081]=16'h6db;
aud[48082]=16'h6f1;
aud[48083]=16'h706;
aud[48084]=16'h71b;
aud[48085]=16'h731;
aud[48086]=16'h746;
aud[48087]=16'h75b;
aud[48088]=16'h770;
aud[48089]=16'h786;
aud[48090]=16'h79b;
aud[48091]=16'h7b0;
aud[48092]=16'h7c6;
aud[48093]=16'h7db;
aud[48094]=16'h7f0;
aud[48095]=16'h805;
aud[48096]=16'h81b;
aud[48097]=16'h830;
aud[48098]=16'h845;
aud[48099]=16'h85b;
aud[48100]=16'h870;
aud[48101]=16'h885;
aud[48102]=16'h89a;
aud[48103]=16'h8b0;
aud[48104]=16'h8c5;
aud[48105]=16'h8da;
aud[48106]=16'h8ef;
aud[48107]=16'h905;
aud[48108]=16'h91a;
aud[48109]=16'h92f;
aud[48110]=16'h944;
aud[48111]=16'h959;
aud[48112]=16'h96f;
aud[48113]=16'h984;
aud[48114]=16'h999;
aud[48115]=16'h9ae;
aud[48116]=16'h9c3;
aud[48117]=16'h9d9;
aud[48118]=16'h9ee;
aud[48119]=16'ha03;
aud[48120]=16'ha18;
aud[48121]=16'ha2d;
aud[48122]=16'ha43;
aud[48123]=16'ha58;
aud[48124]=16'ha6d;
aud[48125]=16'ha82;
aud[48126]=16'ha97;
aud[48127]=16'haac;
aud[48128]=16'hac1;
aud[48129]=16'had7;
aud[48130]=16'haec;
aud[48131]=16'hb01;
aud[48132]=16'hb16;
aud[48133]=16'hb2b;
aud[48134]=16'hb40;
aud[48135]=16'hb55;
aud[48136]=16'hb6a;
aud[48137]=16'hb80;
aud[48138]=16'hb95;
aud[48139]=16'hbaa;
aud[48140]=16'hbbf;
aud[48141]=16'hbd4;
aud[48142]=16'hbe9;
aud[48143]=16'hbfe;
aud[48144]=16'hc13;
aud[48145]=16'hc28;
aud[48146]=16'hc3d;
aud[48147]=16'hc52;
aud[48148]=16'hc67;
aud[48149]=16'hc7c;
aud[48150]=16'hc91;
aud[48151]=16'hca6;
aud[48152]=16'hcbb;
aud[48153]=16'hcd0;
aud[48154]=16'hce5;
aud[48155]=16'hcfa;
aud[48156]=16'hd0f;
aud[48157]=16'hd24;
aud[48158]=16'hd39;
aud[48159]=16'hd4e;
aud[48160]=16'hd63;
aud[48161]=16'hd78;
aud[48162]=16'hd8d;
aud[48163]=16'hda2;
aud[48164]=16'hdb7;
aud[48165]=16'hdcc;
aud[48166]=16'hde1;
aud[48167]=16'hdf6;
aud[48168]=16'he0b;
aud[48169]=16'he20;
aud[48170]=16'he35;
aud[48171]=16'he4a;
aud[48172]=16'he5f;
aud[48173]=16'he74;
aud[48174]=16'he88;
aud[48175]=16'he9d;
aud[48176]=16'heb2;
aud[48177]=16'hec7;
aud[48178]=16'hedc;
aud[48179]=16'hef1;
aud[48180]=16'hf06;
aud[48181]=16'hf1a;
aud[48182]=16'hf2f;
aud[48183]=16'hf44;
aud[48184]=16'hf59;
aud[48185]=16'hf6e;
aud[48186]=16'hf83;
aud[48187]=16'hf97;
aud[48188]=16'hfac;
aud[48189]=16'hfc1;
aud[48190]=16'hfd6;
aud[48191]=16'hfeb;
aud[48192]=16'hfff;
aud[48193]=16'h1014;
aud[48194]=16'h1029;
aud[48195]=16'h103e;
aud[48196]=16'h1052;
aud[48197]=16'h1067;
aud[48198]=16'h107c;
aud[48199]=16'h1090;
aud[48200]=16'h10a5;
aud[48201]=16'h10ba;
aud[48202]=16'h10cf;
aud[48203]=16'h10e3;
aud[48204]=16'h10f8;
aud[48205]=16'h110d;
aud[48206]=16'h1121;
aud[48207]=16'h1136;
aud[48208]=16'h114b;
aud[48209]=16'h115f;
aud[48210]=16'h1174;
aud[48211]=16'h1189;
aud[48212]=16'h119d;
aud[48213]=16'h11b2;
aud[48214]=16'h11c6;
aud[48215]=16'h11db;
aud[48216]=16'h11f0;
aud[48217]=16'h1204;
aud[48218]=16'h1219;
aud[48219]=16'h122d;
aud[48220]=16'h1242;
aud[48221]=16'h1256;
aud[48222]=16'h126b;
aud[48223]=16'h127f;
aud[48224]=16'h1294;
aud[48225]=16'h12a9;
aud[48226]=16'h12bd;
aud[48227]=16'h12d2;
aud[48228]=16'h12e6;
aud[48229]=16'h12fb;
aud[48230]=16'h130f;
aud[48231]=16'h1323;
aud[48232]=16'h1338;
aud[48233]=16'h134c;
aud[48234]=16'h1361;
aud[48235]=16'h1375;
aud[48236]=16'h138a;
aud[48237]=16'h139e;
aud[48238]=16'h13b3;
aud[48239]=16'h13c7;
aud[48240]=16'h13db;
aud[48241]=16'h13f0;
aud[48242]=16'h1404;
aud[48243]=16'h1418;
aud[48244]=16'h142d;
aud[48245]=16'h1441;
aud[48246]=16'h1455;
aud[48247]=16'h146a;
aud[48248]=16'h147e;
aud[48249]=16'h1492;
aud[48250]=16'h14a7;
aud[48251]=16'h14bb;
aud[48252]=16'h14cf;
aud[48253]=16'h14e4;
aud[48254]=16'h14f8;
aud[48255]=16'h150c;
aud[48256]=16'h1520;
aud[48257]=16'h1535;
aud[48258]=16'h1549;
aud[48259]=16'h155d;
aud[48260]=16'h1571;
aud[48261]=16'h1586;
aud[48262]=16'h159a;
aud[48263]=16'h15ae;
aud[48264]=16'h15c2;
aud[48265]=16'h15d6;
aud[48266]=16'h15ea;
aud[48267]=16'h15ff;
aud[48268]=16'h1613;
aud[48269]=16'h1627;
aud[48270]=16'h163b;
aud[48271]=16'h164f;
aud[48272]=16'h1663;
aud[48273]=16'h1677;
aud[48274]=16'h168b;
aud[48275]=16'h169f;
aud[48276]=16'h16b3;
aud[48277]=16'h16c7;
aud[48278]=16'h16db;
aud[48279]=16'h16f0;
aud[48280]=16'h1704;
aud[48281]=16'h1718;
aud[48282]=16'h172c;
aud[48283]=16'h1740;
aud[48284]=16'h1753;
aud[48285]=16'h1767;
aud[48286]=16'h177b;
aud[48287]=16'h178f;
aud[48288]=16'h17a3;
aud[48289]=16'h17b7;
aud[48290]=16'h17cb;
aud[48291]=16'h17df;
aud[48292]=16'h17f3;
aud[48293]=16'h1807;
aud[48294]=16'h181b;
aud[48295]=16'h182f;
aud[48296]=16'h1842;
aud[48297]=16'h1856;
aud[48298]=16'h186a;
aud[48299]=16'h187e;
aud[48300]=16'h1892;
aud[48301]=16'h18a5;
aud[48302]=16'h18b9;
aud[48303]=16'h18cd;
aud[48304]=16'h18e1;
aud[48305]=16'h18f5;
aud[48306]=16'h1908;
aud[48307]=16'h191c;
aud[48308]=16'h1930;
aud[48309]=16'h1943;
aud[48310]=16'h1957;
aud[48311]=16'h196b;
aud[48312]=16'h197f;
aud[48313]=16'h1992;
aud[48314]=16'h19a6;
aud[48315]=16'h19ba;
aud[48316]=16'h19cd;
aud[48317]=16'h19e1;
aud[48318]=16'h19f4;
aud[48319]=16'h1a08;
aud[48320]=16'h1a1c;
aud[48321]=16'h1a2f;
aud[48322]=16'h1a43;
aud[48323]=16'h1a56;
aud[48324]=16'h1a6a;
aud[48325]=16'h1a7d;
aud[48326]=16'h1a91;
aud[48327]=16'h1aa4;
aud[48328]=16'h1ab8;
aud[48329]=16'h1acb;
aud[48330]=16'h1adf;
aud[48331]=16'h1af2;
aud[48332]=16'h1b06;
aud[48333]=16'h1b19;
aud[48334]=16'h1b2d;
aud[48335]=16'h1b40;
aud[48336]=16'h1b53;
aud[48337]=16'h1b67;
aud[48338]=16'h1b7a;
aud[48339]=16'h1b8d;
aud[48340]=16'h1ba1;
aud[48341]=16'h1bb4;
aud[48342]=16'h1bc8;
aud[48343]=16'h1bdb;
aud[48344]=16'h1bee;
aud[48345]=16'h1c01;
aud[48346]=16'h1c15;
aud[48347]=16'h1c28;
aud[48348]=16'h1c3b;
aud[48349]=16'h1c4e;
aud[48350]=16'h1c62;
aud[48351]=16'h1c75;
aud[48352]=16'h1c88;
aud[48353]=16'h1c9b;
aud[48354]=16'h1cae;
aud[48355]=16'h1cc2;
aud[48356]=16'h1cd5;
aud[48357]=16'h1ce8;
aud[48358]=16'h1cfb;
aud[48359]=16'h1d0e;
aud[48360]=16'h1d21;
aud[48361]=16'h1d34;
aud[48362]=16'h1d47;
aud[48363]=16'h1d5b;
aud[48364]=16'h1d6e;
aud[48365]=16'h1d81;
aud[48366]=16'h1d94;
aud[48367]=16'h1da7;
aud[48368]=16'h1dba;
aud[48369]=16'h1dcd;
aud[48370]=16'h1de0;
aud[48371]=16'h1df3;
aud[48372]=16'h1e06;
aud[48373]=16'h1e18;
aud[48374]=16'h1e2b;
aud[48375]=16'h1e3e;
aud[48376]=16'h1e51;
aud[48377]=16'h1e64;
aud[48378]=16'h1e77;
aud[48379]=16'h1e8a;
aud[48380]=16'h1e9d;
aud[48381]=16'h1eaf;
aud[48382]=16'h1ec2;
aud[48383]=16'h1ed5;
aud[48384]=16'h1ee8;
aud[48385]=16'h1efb;
aud[48386]=16'h1f0d;
aud[48387]=16'h1f20;
aud[48388]=16'h1f33;
aud[48389]=16'h1f46;
aud[48390]=16'h1f58;
aud[48391]=16'h1f6b;
aud[48392]=16'h1f7e;
aud[48393]=16'h1f90;
aud[48394]=16'h1fa3;
aud[48395]=16'h1fb6;
aud[48396]=16'h1fc8;
aud[48397]=16'h1fdb;
aud[48398]=16'h1fed;
aud[48399]=16'h2000;
aud[48400]=16'h2013;
aud[48401]=16'h2025;
aud[48402]=16'h2038;
aud[48403]=16'h204a;
aud[48404]=16'h205d;
aud[48405]=16'h206f;
aud[48406]=16'h2082;
aud[48407]=16'h2094;
aud[48408]=16'h20a7;
aud[48409]=16'h20b9;
aud[48410]=16'h20cb;
aud[48411]=16'h20de;
aud[48412]=16'h20f0;
aud[48413]=16'h2103;
aud[48414]=16'h2115;
aud[48415]=16'h2127;
aud[48416]=16'h213a;
aud[48417]=16'h214c;
aud[48418]=16'h215e;
aud[48419]=16'h2171;
aud[48420]=16'h2183;
aud[48421]=16'h2195;
aud[48422]=16'h21a7;
aud[48423]=16'h21ba;
aud[48424]=16'h21cc;
aud[48425]=16'h21de;
aud[48426]=16'h21f0;
aud[48427]=16'h2202;
aud[48428]=16'h2215;
aud[48429]=16'h2227;
aud[48430]=16'h2239;
aud[48431]=16'h224b;
aud[48432]=16'h225d;
aud[48433]=16'h226f;
aud[48434]=16'h2281;
aud[48435]=16'h2293;
aud[48436]=16'h22a5;
aud[48437]=16'h22b7;
aud[48438]=16'h22c9;
aud[48439]=16'h22db;
aud[48440]=16'h22ed;
aud[48441]=16'h22ff;
aud[48442]=16'h2311;
aud[48443]=16'h2323;
aud[48444]=16'h2335;
aud[48445]=16'h2347;
aud[48446]=16'h2359;
aud[48447]=16'h236b;
aud[48448]=16'h237d;
aud[48449]=16'h238e;
aud[48450]=16'h23a0;
aud[48451]=16'h23b2;
aud[48452]=16'h23c4;
aud[48453]=16'h23d6;
aud[48454]=16'h23e7;
aud[48455]=16'h23f9;
aud[48456]=16'h240b;
aud[48457]=16'h241d;
aud[48458]=16'h242e;
aud[48459]=16'h2440;
aud[48460]=16'h2452;
aud[48461]=16'h2463;
aud[48462]=16'h2475;
aud[48463]=16'h2487;
aud[48464]=16'h2498;
aud[48465]=16'h24aa;
aud[48466]=16'h24bb;
aud[48467]=16'h24cd;
aud[48468]=16'h24de;
aud[48469]=16'h24f0;
aud[48470]=16'h2501;
aud[48471]=16'h2513;
aud[48472]=16'h2524;
aud[48473]=16'h2536;
aud[48474]=16'h2547;
aud[48475]=16'h2559;
aud[48476]=16'h256a;
aud[48477]=16'h257c;
aud[48478]=16'h258d;
aud[48479]=16'h259e;
aud[48480]=16'h25b0;
aud[48481]=16'h25c1;
aud[48482]=16'h25d2;
aud[48483]=16'h25e4;
aud[48484]=16'h25f5;
aud[48485]=16'h2606;
aud[48486]=16'h2617;
aud[48487]=16'h2629;
aud[48488]=16'h263a;
aud[48489]=16'h264b;
aud[48490]=16'h265c;
aud[48491]=16'h266d;
aud[48492]=16'h267e;
aud[48493]=16'h2690;
aud[48494]=16'h26a1;
aud[48495]=16'h26b2;
aud[48496]=16'h26c3;
aud[48497]=16'h26d4;
aud[48498]=16'h26e5;
aud[48499]=16'h26f6;
aud[48500]=16'h2707;
aud[48501]=16'h2718;
aud[48502]=16'h2729;
aud[48503]=16'h273a;
aud[48504]=16'h274b;
aud[48505]=16'h275c;
aud[48506]=16'h276d;
aud[48507]=16'h277e;
aud[48508]=16'h278e;
aud[48509]=16'h279f;
aud[48510]=16'h27b0;
aud[48511]=16'h27c1;
aud[48512]=16'h27d2;
aud[48513]=16'h27e2;
aud[48514]=16'h27f3;
aud[48515]=16'h2804;
aud[48516]=16'h2815;
aud[48517]=16'h2825;
aud[48518]=16'h2836;
aud[48519]=16'h2847;
aud[48520]=16'h2857;
aud[48521]=16'h2868;
aud[48522]=16'h2879;
aud[48523]=16'h2889;
aud[48524]=16'h289a;
aud[48525]=16'h28aa;
aud[48526]=16'h28bb;
aud[48527]=16'h28cc;
aud[48528]=16'h28dc;
aud[48529]=16'h28ed;
aud[48530]=16'h28fd;
aud[48531]=16'h290e;
aud[48532]=16'h291e;
aud[48533]=16'h292e;
aud[48534]=16'h293f;
aud[48535]=16'h294f;
aud[48536]=16'h2960;
aud[48537]=16'h2970;
aud[48538]=16'h2980;
aud[48539]=16'h2991;
aud[48540]=16'h29a1;
aud[48541]=16'h29b1;
aud[48542]=16'h29c1;
aud[48543]=16'h29d2;
aud[48544]=16'h29e2;
aud[48545]=16'h29f2;
aud[48546]=16'h2a02;
aud[48547]=16'h2a12;
aud[48548]=16'h2a23;
aud[48549]=16'h2a33;
aud[48550]=16'h2a43;
aud[48551]=16'h2a53;
aud[48552]=16'h2a63;
aud[48553]=16'h2a73;
aud[48554]=16'h2a83;
aud[48555]=16'h2a93;
aud[48556]=16'h2aa3;
aud[48557]=16'h2ab3;
aud[48558]=16'h2ac3;
aud[48559]=16'h2ad3;
aud[48560]=16'h2ae3;
aud[48561]=16'h2af3;
aud[48562]=16'h2b03;
aud[48563]=16'h2b13;
aud[48564]=16'h2b22;
aud[48565]=16'h2b32;
aud[48566]=16'h2b42;
aud[48567]=16'h2b52;
aud[48568]=16'h2b62;
aud[48569]=16'h2b71;
aud[48570]=16'h2b81;
aud[48571]=16'h2b91;
aud[48572]=16'h2ba1;
aud[48573]=16'h2bb0;
aud[48574]=16'h2bc0;
aud[48575]=16'h2bd0;
aud[48576]=16'h2bdf;
aud[48577]=16'h2bef;
aud[48578]=16'h2bfe;
aud[48579]=16'h2c0e;
aud[48580]=16'h2c1e;
aud[48581]=16'h2c2d;
aud[48582]=16'h2c3d;
aud[48583]=16'h2c4c;
aud[48584]=16'h2c5c;
aud[48585]=16'h2c6b;
aud[48586]=16'h2c7a;
aud[48587]=16'h2c8a;
aud[48588]=16'h2c99;
aud[48589]=16'h2ca9;
aud[48590]=16'h2cb8;
aud[48591]=16'h2cc7;
aud[48592]=16'h2cd7;
aud[48593]=16'h2ce6;
aud[48594]=16'h2cf5;
aud[48595]=16'h2d04;
aud[48596]=16'h2d14;
aud[48597]=16'h2d23;
aud[48598]=16'h2d32;
aud[48599]=16'h2d41;
aud[48600]=16'h2d50;
aud[48601]=16'h2d60;
aud[48602]=16'h2d6f;
aud[48603]=16'h2d7e;
aud[48604]=16'h2d8d;
aud[48605]=16'h2d9c;
aud[48606]=16'h2dab;
aud[48607]=16'h2dba;
aud[48608]=16'h2dc9;
aud[48609]=16'h2dd8;
aud[48610]=16'h2de7;
aud[48611]=16'h2df6;
aud[48612]=16'h2e05;
aud[48613]=16'h2e14;
aud[48614]=16'h2e22;
aud[48615]=16'h2e31;
aud[48616]=16'h2e40;
aud[48617]=16'h2e4f;
aud[48618]=16'h2e5e;
aud[48619]=16'h2e6d;
aud[48620]=16'h2e7b;
aud[48621]=16'h2e8a;
aud[48622]=16'h2e99;
aud[48623]=16'h2ea7;
aud[48624]=16'h2eb6;
aud[48625]=16'h2ec5;
aud[48626]=16'h2ed3;
aud[48627]=16'h2ee2;
aud[48628]=16'h2ef1;
aud[48629]=16'h2eff;
aud[48630]=16'h2f0e;
aud[48631]=16'h2f1c;
aud[48632]=16'h2f2b;
aud[48633]=16'h2f39;
aud[48634]=16'h2f48;
aud[48635]=16'h2f56;
aud[48636]=16'h2f65;
aud[48637]=16'h2f73;
aud[48638]=16'h2f81;
aud[48639]=16'h2f90;
aud[48640]=16'h2f9e;
aud[48641]=16'h2fac;
aud[48642]=16'h2fbb;
aud[48643]=16'h2fc9;
aud[48644]=16'h2fd7;
aud[48645]=16'h2fe5;
aud[48646]=16'h2ff4;
aud[48647]=16'h3002;
aud[48648]=16'h3010;
aud[48649]=16'h301e;
aud[48650]=16'h302c;
aud[48651]=16'h303a;
aud[48652]=16'h3048;
aud[48653]=16'h3057;
aud[48654]=16'h3065;
aud[48655]=16'h3073;
aud[48656]=16'h3081;
aud[48657]=16'h308f;
aud[48658]=16'h309d;
aud[48659]=16'h30aa;
aud[48660]=16'h30b8;
aud[48661]=16'h30c6;
aud[48662]=16'h30d4;
aud[48663]=16'h30e2;
aud[48664]=16'h30f0;
aud[48665]=16'h30fe;
aud[48666]=16'h310b;
aud[48667]=16'h3119;
aud[48668]=16'h3127;
aud[48669]=16'h3135;
aud[48670]=16'h3142;
aud[48671]=16'h3150;
aud[48672]=16'h315e;
aud[48673]=16'h316b;
aud[48674]=16'h3179;
aud[48675]=16'h3187;
aud[48676]=16'h3194;
aud[48677]=16'h31a2;
aud[48678]=16'h31af;
aud[48679]=16'h31bd;
aud[48680]=16'h31ca;
aud[48681]=16'h31d8;
aud[48682]=16'h31e5;
aud[48683]=16'h31f3;
aud[48684]=16'h3200;
aud[48685]=16'h320d;
aud[48686]=16'h321b;
aud[48687]=16'h3228;
aud[48688]=16'h3235;
aud[48689]=16'h3243;
aud[48690]=16'h3250;
aud[48691]=16'h325d;
aud[48692]=16'h326a;
aud[48693]=16'h3278;
aud[48694]=16'h3285;
aud[48695]=16'h3292;
aud[48696]=16'h329f;
aud[48697]=16'h32ac;
aud[48698]=16'h32b9;
aud[48699]=16'h32c6;
aud[48700]=16'h32d3;
aud[48701]=16'h32e0;
aud[48702]=16'h32ed;
aud[48703]=16'h32fa;
aud[48704]=16'h3307;
aud[48705]=16'h3314;
aud[48706]=16'h3321;
aud[48707]=16'h332e;
aud[48708]=16'h333b;
aud[48709]=16'h3348;
aud[48710]=16'h3355;
aud[48711]=16'h3361;
aud[48712]=16'h336e;
aud[48713]=16'h337b;
aud[48714]=16'h3388;
aud[48715]=16'h3394;
aud[48716]=16'h33a1;
aud[48717]=16'h33ae;
aud[48718]=16'h33ba;
aud[48719]=16'h33c7;
aud[48720]=16'h33d4;
aud[48721]=16'h33e0;
aud[48722]=16'h33ed;
aud[48723]=16'h33f9;
aud[48724]=16'h3406;
aud[48725]=16'h3412;
aud[48726]=16'h341f;
aud[48727]=16'h342b;
aud[48728]=16'h3437;
aud[48729]=16'h3444;
aud[48730]=16'h3450;
aud[48731]=16'h345d;
aud[48732]=16'h3469;
aud[48733]=16'h3475;
aud[48734]=16'h3481;
aud[48735]=16'h348e;
aud[48736]=16'h349a;
aud[48737]=16'h34a6;
aud[48738]=16'h34b2;
aud[48739]=16'h34be;
aud[48740]=16'h34cb;
aud[48741]=16'h34d7;
aud[48742]=16'h34e3;
aud[48743]=16'h34ef;
aud[48744]=16'h34fb;
aud[48745]=16'h3507;
aud[48746]=16'h3513;
aud[48747]=16'h351f;
aud[48748]=16'h352b;
aud[48749]=16'h3537;
aud[48750]=16'h3543;
aud[48751]=16'h354f;
aud[48752]=16'h355a;
aud[48753]=16'h3566;
aud[48754]=16'h3572;
aud[48755]=16'h357e;
aud[48756]=16'h358a;
aud[48757]=16'h3595;
aud[48758]=16'h35a1;
aud[48759]=16'h35ad;
aud[48760]=16'h35b8;
aud[48761]=16'h35c4;
aud[48762]=16'h35d0;
aud[48763]=16'h35db;
aud[48764]=16'h35e7;
aud[48765]=16'h35f2;
aud[48766]=16'h35fe;
aud[48767]=16'h3609;
aud[48768]=16'h3615;
aud[48769]=16'h3620;
aud[48770]=16'h362c;
aud[48771]=16'h3637;
aud[48772]=16'h3643;
aud[48773]=16'h364e;
aud[48774]=16'h3659;
aud[48775]=16'h3665;
aud[48776]=16'h3670;
aud[48777]=16'h367b;
aud[48778]=16'h3686;
aud[48779]=16'h3692;
aud[48780]=16'h369d;
aud[48781]=16'h36a8;
aud[48782]=16'h36b3;
aud[48783]=16'h36be;
aud[48784]=16'h36c9;
aud[48785]=16'h36d4;
aud[48786]=16'h36e0;
aud[48787]=16'h36eb;
aud[48788]=16'h36f6;
aud[48789]=16'h3701;
aud[48790]=16'h370b;
aud[48791]=16'h3716;
aud[48792]=16'h3721;
aud[48793]=16'h372c;
aud[48794]=16'h3737;
aud[48795]=16'h3742;
aud[48796]=16'h374d;
aud[48797]=16'h3757;
aud[48798]=16'h3762;
aud[48799]=16'h376d;
aud[48800]=16'h3778;
aud[48801]=16'h3782;
aud[48802]=16'h378d;
aud[48803]=16'h3798;
aud[48804]=16'h37a2;
aud[48805]=16'h37ad;
aud[48806]=16'h37b7;
aud[48807]=16'h37c2;
aud[48808]=16'h37cc;
aud[48809]=16'h37d7;
aud[48810]=16'h37e1;
aud[48811]=16'h37ec;
aud[48812]=16'h37f6;
aud[48813]=16'h3801;
aud[48814]=16'h380b;
aud[48815]=16'h3815;
aud[48816]=16'h3820;
aud[48817]=16'h382a;
aud[48818]=16'h3834;
aud[48819]=16'h383f;
aud[48820]=16'h3849;
aud[48821]=16'h3853;
aud[48822]=16'h385d;
aud[48823]=16'h3867;
aud[48824]=16'h3871;
aud[48825]=16'h387b;
aud[48826]=16'h3886;
aud[48827]=16'h3890;
aud[48828]=16'h389a;
aud[48829]=16'h38a4;
aud[48830]=16'h38ae;
aud[48831]=16'h38b8;
aud[48832]=16'h38c1;
aud[48833]=16'h38cb;
aud[48834]=16'h38d5;
aud[48835]=16'h38df;
aud[48836]=16'h38e9;
aud[48837]=16'h38f3;
aud[48838]=16'h38fd;
aud[48839]=16'h3906;
aud[48840]=16'h3910;
aud[48841]=16'h391a;
aud[48842]=16'h3923;
aud[48843]=16'h392d;
aud[48844]=16'h3937;
aud[48845]=16'h3940;
aud[48846]=16'h394a;
aud[48847]=16'h3953;
aud[48848]=16'h395d;
aud[48849]=16'h3966;
aud[48850]=16'h3970;
aud[48851]=16'h3979;
aud[48852]=16'h3983;
aud[48853]=16'h398c;
aud[48854]=16'h3995;
aud[48855]=16'h399f;
aud[48856]=16'h39a8;
aud[48857]=16'h39b1;
aud[48858]=16'h39bb;
aud[48859]=16'h39c4;
aud[48860]=16'h39cd;
aud[48861]=16'h39d6;
aud[48862]=16'h39e0;
aud[48863]=16'h39e9;
aud[48864]=16'h39f2;
aud[48865]=16'h39fb;
aud[48866]=16'h3a04;
aud[48867]=16'h3a0d;
aud[48868]=16'h3a16;
aud[48869]=16'h3a1f;
aud[48870]=16'h3a28;
aud[48871]=16'h3a31;
aud[48872]=16'h3a3a;
aud[48873]=16'h3a43;
aud[48874]=16'h3a4c;
aud[48875]=16'h3a54;
aud[48876]=16'h3a5d;
aud[48877]=16'h3a66;
aud[48878]=16'h3a6f;
aud[48879]=16'h3a78;
aud[48880]=16'h3a80;
aud[48881]=16'h3a89;
aud[48882]=16'h3a92;
aud[48883]=16'h3a9a;
aud[48884]=16'h3aa3;
aud[48885]=16'h3aab;
aud[48886]=16'h3ab4;
aud[48887]=16'h3abc;
aud[48888]=16'h3ac5;
aud[48889]=16'h3acd;
aud[48890]=16'h3ad6;
aud[48891]=16'h3ade;
aud[48892]=16'h3ae7;
aud[48893]=16'h3aef;
aud[48894]=16'h3af7;
aud[48895]=16'h3b00;
aud[48896]=16'h3b08;
aud[48897]=16'h3b10;
aud[48898]=16'h3b19;
aud[48899]=16'h3b21;
aud[48900]=16'h3b29;
aud[48901]=16'h3b31;
aud[48902]=16'h3b39;
aud[48903]=16'h3b41;
aud[48904]=16'h3b4a;
aud[48905]=16'h3b52;
aud[48906]=16'h3b5a;
aud[48907]=16'h3b62;
aud[48908]=16'h3b6a;
aud[48909]=16'h3b72;
aud[48910]=16'h3b7a;
aud[48911]=16'h3b81;
aud[48912]=16'h3b89;
aud[48913]=16'h3b91;
aud[48914]=16'h3b99;
aud[48915]=16'h3ba1;
aud[48916]=16'h3ba9;
aud[48917]=16'h3bb0;
aud[48918]=16'h3bb8;
aud[48919]=16'h3bc0;
aud[48920]=16'h3bc7;
aud[48921]=16'h3bcf;
aud[48922]=16'h3bd7;
aud[48923]=16'h3bde;
aud[48924]=16'h3be6;
aud[48925]=16'h3bed;
aud[48926]=16'h3bf5;
aud[48927]=16'h3bfc;
aud[48928]=16'h3c04;
aud[48929]=16'h3c0b;
aud[48930]=16'h3c13;
aud[48931]=16'h3c1a;
aud[48932]=16'h3c21;
aud[48933]=16'h3c29;
aud[48934]=16'h3c30;
aud[48935]=16'h3c37;
aud[48936]=16'h3c3f;
aud[48937]=16'h3c46;
aud[48938]=16'h3c4d;
aud[48939]=16'h3c54;
aud[48940]=16'h3c5b;
aud[48941]=16'h3c63;
aud[48942]=16'h3c6a;
aud[48943]=16'h3c71;
aud[48944]=16'h3c78;
aud[48945]=16'h3c7f;
aud[48946]=16'h3c86;
aud[48947]=16'h3c8d;
aud[48948]=16'h3c94;
aud[48949]=16'h3c9b;
aud[48950]=16'h3ca1;
aud[48951]=16'h3ca8;
aud[48952]=16'h3caf;
aud[48953]=16'h3cb6;
aud[48954]=16'h3cbd;
aud[48955]=16'h3cc3;
aud[48956]=16'h3cca;
aud[48957]=16'h3cd1;
aud[48958]=16'h3cd7;
aud[48959]=16'h3cde;
aud[48960]=16'h3ce5;
aud[48961]=16'h3ceb;
aud[48962]=16'h3cf2;
aud[48963]=16'h3cf8;
aud[48964]=16'h3cff;
aud[48965]=16'h3d05;
aud[48966]=16'h3d0c;
aud[48967]=16'h3d12;
aud[48968]=16'h3d19;
aud[48969]=16'h3d1f;
aud[48970]=16'h3d25;
aud[48971]=16'h3d2c;
aud[48972]=16'h3d32;
aud[48973]=16'h3d38;
aud[48974]=16'h3d3f;
aud[48975]=16'h3d45;
aud[48976]=16'h3d4b;
aud[48977]=16'h3d51;
aud[48978]=16'h3d57;
aud[48979]=16'h3d5d;
aud[48980]=16'h3d63;
aud[48981]=16'h3d69;
aud[48982]=16'h3d6f;
aud[48983]=16'h3d75;
aud[48984]=16'h3d7b;
aud[48985]=16'h3d81;
aud[48986]=16'h3d87;
aud[48987]=16'h3d8d;
aud[48988]=16'h3d93;
aud[48989]=16'h3d99;
aud[48990]=16'h3d9f;
aud[48991]=16'h3da4;
aud[48992]=16'h3daa;
aud[48993]=16'h3db0;
aud[48994]=16'h3db6;
aud[48995]=16'h3dbb;
aud[48996]=16'h3dc1;
aud[48997]=16'h3dc7;
aud[48998]=16'h3dcc;
aud[48999]=16'h3dd2;
aud[49000]=16'h3dd7;
aud[49001]=16'h3ddd;
aud[49002]=16'h3de2;
aud[49003]=16'h3de8;
aud[49004]=16'h3ded;
aud[49005]=16'h3df3;
aud[49006]=16'h3df8;
aud[49007]=16'h3dfd;
aud[49008]=16'h3e03;
aud[49009]=16'h3e08;
aud[49010]=16'h3e0d;
aud[49011]=16'h3e12;
aud[49012]=16'h3e18;
aud[49013]=16'h3e1d;
aud[49014]=16'h3e22;
aud[49015]=16'h3e27;
aud[49016]=16'h3e2c;
aud[49017]=16'h3e31;
aud[49018]=16'h3e36;
aud[49019]=16'h3e3b;
aud[49020]=16'h3e40;
aud[49021]=16'h3e45;
aud[49022]=16'h3e4a;
aud[49023]=16'h3e4f;
aud[49024]=16'h3e54;
aud[49025]=16'h3e59;
aud[49026]=16'h3e5e;
aud[49027]=16'h3e62;
aud[49028]=16'h3e67;
aud[49029]=16'h3e6c;
aud[49030]=16'h3e71;
aud[49031]=16'h3e75;
aud[49032]=16'h3e7a;
aud[49033]=16'h3e7f;
aud[49034]=16'h3e83;
aud[49035]=16'h3e88;
aud[49036]=16'h3e8c;
aud[49037]=16'h3e91;
aud[49038]=16'h3e95;
aud[49039]=16'h3e9a;
aud[49040]=16'h3e9e;
aud[49041]=16'h3ea3;
aud[49042]=16'h3ea7;
aud[49043]=16'h3eac;
aud[49044]=16'h3eb0;
aud[49045]=16'h3eb4;
aud[49046]=16'h3eb9;
aud[49047]=16'h3ebd;
aud[49048]=16'h3ec1;
aud[49049]=16'h3ec5;
aud[49050]=16'h3ec9;
aud[49051]=16'h3ecd;
aud[49052]=16'h3ed2;
aud[49053]=16'h3ed6;
aud[49054]=16'h3eda;
aud[49055]=16'h3ede;
aud[49056]=16'h3ee2;
aud[49057]=16'h3ee6;
aud[49058]=16'h3eea;
aud[49059]=16'h3eee;
aud[49060]=16'h3ef2;
aud[49061]=16'h3ef5;
aud[49062]=16'h3ef9;
aud[49063]=16'h3efd;
aud[49064]=16'h3f01;
aud[49065]=16'h3f05;
aud[49066]=16'h3f08;
aud[49067]=16'h3f0c;
aud[49068]=16'h3f10;
aud[49069]=16'h3f13;
aud[49070]=16'h3f17;
aud[49071]=16'h3f1b;
aud[49072]=16'h3f1e;
aud[49073]=16'h3f22;
aud[49074]=16'h3f25;
aud[49075]=16'h3f29;
aud[49076]=16'h3f2c;
aud[49077]=16'h3f30;
aud[49078]=16'h3f33;
aud[49079]=16'h3f36;
aud[49080]=16'h3f3a;
aud[49081]=16'h3f3d;
aud[49082]=16'h3f40;
aud[49083]=16'h3f43;
aud[49084]=16'h3f47;
aud[49085]=16'h3f4a;
aud[49086]=16'h3f4d;
aud[49087]=16'h3f50;
aud[49088]=16'h3f53;
aud[49089]=16'h3f56;
aud[49090]=16'h3f5a;
aud[49091]=16'h3f5d;
aud[49092]=16'h3f60;
aud[49093]=16'h3f63;
aud[49094]=16'h3f65;
aud[49095]=16'h3f68;
aud[49096]=16'h3f6b;
aud[49097]=16'h3f6e;
aud[49098]=16'h3f71;
aud[49099]=16'h3f74;
aud[49100]=16'h3f77;
aud[49101]=16'h3f79;
aud[49102]=16'h3f7c;
aud[49103]=16'h3f7f;
aud[49104]=16'h3f81;
aud[49105]=16'h3f84;
aud[49106]=16'h3f87;
aud[49107]=16'h3f89;
aud[49108]=16'h3f8c;
aud[49109]=16'h3f8e;
aud[49110]=16'h3f91;
aud[49111]=16'h3f93;
aud[49112]=16'h3f96;
aud[49113]=16'h3f98;
aud[49114]=16'h3f9b;
aud[49115]=16'h3f9d;
aud[49116]=16'h3f9f;
aud[49117]=16'h3fa2;
aud[49118]=16'h3fa4;
aud[49119]=16'h3fa6;
aud[49120]=16'h3fa8;
aud[49121]=16'h3fab;
aud[49122]=16'h3fad;
aud[49123]=16'h3faf;
aud[49124]=16'h3fb1;
aud[49125]=16'h3fb3;
aud[49126]=16'h3fb5;
aud[49127]=16'h3fb7;
aud[49128]=16'h3fb9;
aud[49129]=16'h3fbb;
aud[49130]=16'h3fbd;
aud[49131]=16'h3fbf;
aud[49132]=16'h3fc1;
aud[49133]=16'h3fc3;
aud[49134]=16'h3fc5;
aud[49135]=16'h3fc7;
aud[49136]=16'h3fc8;
aud[49137]=16'h3fca;
aud[49138]=16'h3fcc;
aud[49139]=16'h3fcd;
aud[49140]=16'h3fcf;
aud[49141]=16'h3fd1;
aud[49142]=16'h3fd2;
aud[49143]=16'h3fd4;
aud[49144]=16'h3fd6;
aud[49145]=16'h3fd7;
aud[49146]=16'h3fd9;
aud[49147]=16'h3fda;
aud[49148]=16'h3fdc;
aud[49149]=16'h3fdd;
aud[49150]=16'h3fde;
aud[49151]=16'h3fe0;
aud[49152]=16'h3fe1;
aud[49153]=16'h3fe2;
aud[49154]=16'h3fe4;
aud[49155]=16'h3fe5;
aud[49156]=16'h3fe6;
aud[49157]=16'h3fe7;
aud[49158]=16'h3fe8;
aud[49159]=16'h3fea;
aud[49160]=16'h3feb;
aud[49161]=16'h3fec;
aud[49162]=16'h3fed;
aud[49163]=16'h3fee;
aud[49164]=16'h3fef;
aud[49165]=16'h3ff0;
aud[49166]=16'h3ff1;
aud[49167]=16'h3ff2;
aud[49168]=16'h3ff3;
aud[49169]=16'h3ff3;
aud[49170]=16'h3ff4;
aud[49171]=16'h3ff5;
aud[49172]=16'h3ff6;
aud[49173]=16'h3ff7;
aud[49174]=16'h3ff7;
aud[49175]=16'h3ff8;
aud[49176]=16'h3ff9;
aud[49177]=16'h3ff9;
aud[49178]=16'h3ffa;
aud[49179]=16'h3ffa;
aud[49180]=16'h3ffb;
aud[49181]=16'h3ffb;
aud[49182]=16'h3ffc;
aud[49183]=16'h3ffc;
aud[49184]=16'h3ffd;
aud[49185]=16'h3ffd;
aud[49186]=16'h3ffe;
aud[49187]=16'h3ffe;
aud[49188]=16'h3ffe;
aud[49189]=16'h3fff;
aud[49190]=16'h3fff;
aud[49191]=16'h3fff;
aud[49192]=16'h3fff;
aud[49193]=16'h3fff;
aud[49194]=16'h4000;
aud[49195]=16'h4000;
aud[49196]=16'h4000;
aud[49197]=16'h4000;
aud[49198]=16'h4000;
aud[49199]=16'h4000;
aud[49200]=16'h4000;
aud[49201]=16'h4000;
aud[49202]=16'h4000;
aud[49203]=16'h4000;
aud[49204]=16'h4000;
aud[49205]=16'h3fff;
aud[49206]=16'h3fff;
aud[49207]=16'h3fff;
aud[49208]=16'h3fff;
aud[49209]=16'h3fff;
aud[49210]=16'h3ffe;
aud[49211]=16'h3ffe;
aud[49212]=16'h3ffe;
aud[49213]=16'h3ffd;
aud[49214]=16'h3ffd;
aud[49215]=16'h3ffc;
aud[49216]=16'h3ffc;
aud[49217]=16'h3ffb;
aud[49218]=16'h3ffb;
aud[49219]=16'h3ffa;
aud[49220]=16'h3ffa;
aud[49221]=16'h3ff9;
aud[49222]=16'h3ff9;
aud[49223]=16'h3ff8;
aud[49224]=16'h3ff7;
aud[49225]=16'h3ff7;
aud[49226]=16'h3ff6;
aud[49227]=16'h3ff5;
aud[49228]=16'h3ff4;
aud[49229]=16'h3ff3;
aud[49230]=16'h3ff3;
aud[49231]=16'h3ff2;
aud[49232]=16'h3ff1;
aud[49233]=16'h3ff0;
aud[49234]=16'h3fef;
aud[49235]=16'h3fee;
aud[49236]=16'h3fed;
aud[49237]=16'h3fec;
aud[49238]=16'h3feb;
aud[49239]=16'h3fea;
aud[49240]=16'h3fe8;
aud[49241]=16'h3fe7;
aud[49242]=16'h3fe6;
aud[49243]=16'h3fe5;
aud[49244]=16'h3fe4;
aud[49245]=16'h3fe2;
aud[49246]=16'h3fe1;
aud[49247]=16'h3fe0;
aud[49248]=16'h3fde;
aud[49249]=16'h3fdd;
aud[49250]=16'h3fdc;
aud[49251]=16'h3fda;
aud[49252]=16'h3fd9;
aud[49253]=16'h3fd7;
aud[49254]=16'h3fd6;
aud[49255]=16'h3fd4;
aud[49256]=16'h3fd2;
aud[49257]=16'h3fd1;
aud[49258]=16'h3fcf;
aud[49259]=16'h3fcd;
aud[49260]=16'h3fcc;
aud[49261]=16'h3fca;
aud[49262]=16'h3fc8;
aud[49263]=16'h3fc7;
aud[49264]=16'h3fc5;
aud[49265]=16'h3fc3;
aud[49266]=16'h3fc1;
aud[49267]=16'h3fbf;
aud[49268]=16'h3fbd;
aud[49269]=16'h3fbb;
aud[49270]=16'h3fb9;
aud[49271]=16'h3fb7;
aud[49272]=16'h3fb5;
aud[49273]=16'h3fb3;
aud[49274]=16'h3fb1;
aud[49275]=16'h3faf;
aud[49276]=16'h3fad;
aud[49277]=16'h3fab;
aud[49278]=16'h3fa8;
aud[49279]=16'h3fa6;
aud[49280]=16'h3fa4;
aud[49281]=16'h3fa2;
aud[49282]=16'h3f9f;
aud[49283]=16'h3f9d;
aud[49284]=16'h3f9b;
aud[49285]=16'h3f98;
aud[49286]=16'h3f96;
aud[49287]=16'h3f93;
aud[49288]=16'h3f91;
aud[49289]=16'h3f8e;
aud[49290]=16'h3f8c;
aud[49291]=16'h3f89;
aud[49292]=16'h3f87;
aud[49293]=16'h3f84;
aud[49294]=16'h3f81;
aud[49295]=16'h3f7f;
aud[49296]=16'h3f7c;
aud[49297]=16'h3f79;
aud[49298]=16'h3f77;
aud[49299]=16'h3f74;
aud[49300]=16'h3f71;
aud[49301]=16'h3f6e;
aud[49302]=16'h3f6b;
aud[49303]=16'h3f68;
aud[49304]=16'h3f65;
aud[49305]=16'h3f63;
aud[49306]=16'h3f60;
aud[49307]=16'h3f5d;
aud[49308]=16'h3f5a;
aud[49309]=16'h3f56;
aud[49310]=16'h3f53;
aud[49311]=16'h3f50;
aud[49312]=16'h3f4d;
aud[49313]=16'h3f4a;
aud[49314]=16'h3f47;
aud[49315]=16'h3f43;
aud[49316]=16'h3f40;
aud[49317]=16'h3f3d;
aud[49318]=16'h3f3a;
aud[49319]=16'h3f36;
aud[49320]=16'h3f33;
aud[49321]=16'h3f30;
aud[49322]=16'h3f2c;
aud[49323]=16'h3f29;
aud[49324]=16'h3f25;
aud[49325]=16'h3f22;
aud[49326]=16'h3f1e;
aud[49327]=16'h3f1b;
aud[49328]=16'h3f17;
aud[49329]=16'h3f13;
aud[49330]=16'h3f10;
aud[49331]=16'h3f0c;
aud[49332]=16'h3f08;
aud[49333]=16'h3f05;
aud[49334]=16'h3f01;
aud[49335]=16'h3efd;
aud[49336]=16'h3ef9;
aud[49337]=16'h3ef5;
aud[49338]=16'h3ef2;
aud[49339]=16'h3eee;
aud[49340]=16'h3eea;
aud[49341]=16'h3ee6;
aud[49342]=16'h3ee2;
aud[49343]=16'h3ede;
aud[49344]=16'h3eda;
aud[49345]=16'h3ed6;
aud[49346]=16'h3ed2;
aud[49347]=16'h3ecd;
aud[49348]=16'h3ec9;
aud[49349]=16'h3ec5;
aud[49350]=16'h3ec1;
aud[49351]=16'h3ebd;
aud[49352]=16'h3eb9;
aud[49353]=16'h3eb4;
aud[49354]=16'h3eb0;
aud[49355]=16'h3eac;
aud[49356]=16'h3ea7;
aud[49357]=16'h3ea3;
aud[49358]=16'h3e9e;
aud[49359]=16'h3e9a;
aud[49360]=16'h3e95;
aud[49361]=16'h3e91;
aud[49362]=16'h3e8c;
aud[49363]=16'h3e88;
aud[49364]=16'h3e83;
aud[49365]=16'h3e7f;
aud[49366]=16'h3e7a;
aud[49367]=16'h3e75;
aud[49368]=16'h3e71;
aud[49369]=16'h3e6c;
aud[49370]=16'h3e67;
aud[49371]=16'h3e62;
aud[49372]=16'h3e5e;
aud[49373]=16'h3e59;
aud[49374]=16'h3e54;
aud[49375]=16'h3e4f;
aud[49376]=16'h3e4a;
aud[49377]=16'h3e45;
aud[49378]=16'h3e40;
aud[49379]=16'h3e3b;
aud[49380]=16'h3e36;
aud[49381]=16'h3e31;
aud[49382]=16'h3e2c;
aud[49383]=16'h3e27;
aud[49384]=16'h3e22;
aud[49385]=16'h3e1d;
aud[49386]=16'h3e18;
aud[49387]=16'h3e12;
aud[49388]=16'h3e0d;
aud[49389]=16'h3e08;
aud[49390]=16'h3e03;
aud[49391]=16'h3dfd;
aud[49392]=16'h3df8;
aud[49393]=16'h3df3;
aud[49394]=16'h3ded;
aud[49395]=16'h3de8;
aud[49396]=16'h3de2;
aud[49397]=16'h3ddd;
aud[49398]=16'h3dd7;
aud[49399]=16'h3dd2;
aud[49400]=16'h3dcc;
aud[49401]=16'h3dc7;
aud[49402]=16'h3dc1;
aud[49403]=16'h3dbb;
aud[49404]=16'h3db6;
aud[49405]=16'h3db0;
aud[49406]=16'h3daa;
aud[49407]=16'h3da4;
aud[49408]=16'h3d9f;
aud[49409]=16'h3d99;
aud[49410]=16'h3d93;
aud[49411]=16'h3d8d;
aud[49412]=16'h3d87;
aud[49413]=16'h3d81;
aud[49414]=16'h3d7b;
aud[49415]=16'h3d75;
aud[49416]=16'h3d6f;
aud[49417]=16'h3d69;
aud[49418]=16'h3d63;
aud[49419]=16'h3d5d;
aud[49420]=16'h3d57;
aud[49421]=16'h3d51;
aud[49422]=16'h3d4b;
aud[49423]=16'h3d45;
aud[49424]=16'h3d3f;
aud[49425]=16'h3d38;
aud[49426]=16'h3d32;
aud[49427]=16'h3d2c;
aud[49428]=16'h3d25;
aud[49429]=16'h3d1f;
aud[49430]=16'h3d19;
aud[49431]=16'h3d12;
aud[49432]=16'h3d0c;
aud[49433]=16'h3d05;
aud[49434]=16'h3cff;
aud[49435]=16'h3cf8;
aud[49436]=16'h3cf2;
aud[49437]=16'h3ceb;
aud[49438]=16'h3ce5;
aud[49439]=16'h3cde;
aud[49440]=16'h3cd7;
aud[49441]=16'h3cd1;
aud[49442]=16'h3cca;
aud[49443]=16'h3cc3;
aud[49444]=16'h3cbd;
aud[49445]=16'h3cb6;
aud[49446]=16'h3caf;
aud[49447]=16'h3ca8;
aud[49448]=16'h3ca1;
aud[49449]=16'h3c9b;
aud[49450]=16'h3c94;
aud[49451]=16'h3c8d;
aud[49452]=16'h3c86;
aud[49453]=16'h3c7f;
aud[49454]=16'h3c78;
aud[49455]=16'h3c71;
aud[49456]=16'h3c6a;
aud[49457]=16'h3c63;
aud[49458]=16'h3c5b;
aud[49459]=16'h3c54;
aud[49460]=16'h3c4d;
aud[49461]=16'h3c46;
aud[49462]=16'h3c3f;
aud[49463]=16'h3c37;
aud[49464]=16'h3c30;
aud[49465]=16'h3c29;
aud[49466]=16'h3c21;
aud[49467]=16'h3c1a;
aud[49468]=16'h3c13;
aud[49469]=16'h3c0b;
aud[49470]=16'h3c04;
aud[49471]=16'h3bfc;
aud[49472]=16'h3bf5;
aud[49473]=16'h3bed;
aud[49474]=16'h3be6;
aud[49475]=16'h3bde;
aud[49476]=16'h3bd7;
aud[49477]=16'h3bcf;
aud[49478]=16'h3bc7;
aud[49479]=16'h3bc0;
aud[49480]=16'h3bb8;
aud[49481]=16'h3bb0;
aud[49482]=16'h3ba9;
aud[49483]=16'h3ba1;
aud[49484]=16'h3b99;
aud[49485]=16'h3b91;
aud[49486]=16'h3b89;
aud[49487]=16'h3b81;
aud[49488]=16'h3b7a;
aud[49489]=16'h3b72;
aud[49490]=16'h3b6a;
aud[49491]=16'h3b62;
aud[49492]=16'h3b5a;
aud[49493]=16'h3b52;
aud[49494]=16'h3b4a;
aud[49495]=16'h3b41;
aud[49496]=16'h3b39;
aud[49497]=16'h3b31;
aud[49498]=16'h3b29;
aud[49499]=16'h3b21;
aud[49500]=16'h3b19;
aud[49501]=16'h3b10;
aud[49502]=16'h3b08;
aud[49503]=16'h3b00;
aud[49504]=16'h3af7;
aud[49505]=16'h3aef;
aud[49506]=16'h3ae7;
aud[49507]=16'h3ade;
aud[49508]=16'h3ad6;
aud[49509]=16'h3acd;
aud[49510]=16'h3ac5;
aud[49511]=16'h3abc;
aud[49512]=16'h3ab4;
aud[49513]=16'h3aab;
aud[49514]=16'h3aa3;
aud[49515]=16'h3a9a;
aud[49516]=16'h3a92;
aud[49517]=16'h3a89;
aud[49518]=16'h3a80;
aud[49519]=16'h3a78;
aud[49520]=16'h3a6f;
aud[49521]=16'h3a66;
aud[49522]=16'h3a5d;
aud[49523]=16'h3a54;
aud[49524]=16'h3a4c;
aud[49525]=16'h3a43;
aud[49526]=16'h3a3a;
aud[49527]=16'h3a31;
aud[49528]=16'h3a28;
aud[49529]=16'h3a1f;
aud[49530]=16'h3a16;
aud[49531]=16'h3a0d;
aud[49532]=16'h3a04;
aud[49533]=16'h39fb;
aud[49534]=16'h39f2;
aud[49535]=16'h39e9;
aud[49536]=16'h39e0;
aud[49537]=16'h39d6;
aud[49538]=16'h39cd;
aud[49539]=16'h39c4;
aud[49540]=16'h39bb;
aud[49541]=16'h39b1;
aud[49542]=16'h39a8;
aud[49543]=16'h399f;
aud[49544]=16'h3995;
aud[49545]=16'h398c;
aud[49546]=16'h3983;
aud[49547]=16'h3979;
aud[49548]=16'h3970;
aud[49549]=16'h3966;
aud[49550]=16'h395d;
aud[49551]=16'h3953;
aud[49552]=16'h394a;
aud[49553]=16'h3940;
aud[49554]=16'h3937;
aud[49555]=16'h392d;
aud[49556]=16'h3923;
aud[49557]=16'h391a;
aud[49558]=16'h3910;
aud[49559]=16'h3906;
aud[49560]=16'h38fd;
aud[49561]=16'h38f3;
aud[49562]=16'h38e9;
aud[49563]=16'h38df;
aud[49564]=16'h38d5;
aud[49565]=16'h38cb;
aud[49566]=16'h38c1;
aud[49567]=16'h38b8;
aud[49568]=16'h38ae;
aud[49569]=16'h38a4;
aud[49570]=16'h389a;
aud[49571]=16'h3890;
aud[49572]=16'h3886;
aud[49573]=16'h387b;
aud[49574]=16'h3871;
aud[49575]=16'h3867;
aud[49576]=16'h385d;
aud[49577]=16'h3853;
aud[49578]=16'h3849;
aud[49579]=16'h383f;
aud[49580]=16'h3834;
aud[49581]=16'h382a;
aud[49582]=16'h3820;
aud[49583]=16'h3815;
aud[49584]=16'h380b;
aud[49585]=16'h3801;
aud[49586]=16'h37f6;
aud[49587]=16'h37ec;
aud[49588]=16'h37e1;
aud[49589]=16'h37d7;
aud[49590]=16'h37cc;
aud[49591]=16'h37c2;
aud[49592]=16'h37b7;
aud[49593]=16'h37ad;
aud[49594]=16'h37a2;
aud[49595]=16'h3798;
aud[49596]=16'h378d;
aud[49597]=16'h3782;
aud[49598]=16'h3778;
aud[49599]=16'h376d;
aud[49600]=16'h3762;
aud[49601]=16'h3757;
aud[49602]=16'h374d;
aud[49603]=16'h3742;
aud[49604]=16'h3737;
aud[49605]=16'h372c;
aud[49606]=16'h3721;
aud[49607]=16'h3716;
aud[49608]=16'h370b;
aud[49609]=16'h3701;
aud[49610]=16'h36f6;
aud[49611]=16'h36eb;
aud[49612]=16'h36e0;
aud[49613]=16'h36d4;
aud[49614]=16'h36c9;
aud[49615]=16'h36be;
aud[49616]=16'h36b3;
aud[49617]=16'h36a8;
aud[49618]=16'h369d;
aud[49619]=16'h3692;
aud[49620]=16'h3686;
aud[49621]=16'h367b;
aud[49622]=16'h3670;
aud[49623]=16'h3665;
aud[49624]=16'h3659;
aud[49625]=16'h364e;
aud[49626]=16'h3643;
aud[49627]=16'h3637;
aud[49628]=16'h362c;
aud[49629]=16'h3620;
aud[49630]=16'h3615;
aud[49631]=16'h3609;
aud[49632]=16'h35fe;
aud[49633]=16'h35f2;
aud[49634]=16'h35e7;
aud[49635]=16'h35db;
aud[49636]=16'h35d0;
aud[49637]=16'h35c4;
aud[49638]=16'h35b8;
aud[49639]=16'h35ad;
aud[49640]=16'h35a1;
aud[49641]=16'h3595;
aud[49642]=16'h358a;
aud[49643]=16'h357e;
aud[49644]=16'h3572;
aud[49645]=16'h3566;
aud[49646]=16'h355a;
aud[49647]=16'h354f;
aud[49648]=16'h3543;
aud[49649]=16'h3537;
aud[49650]=16'h352b;
aud[49651]=16'h351f;
aud[49652]=16'h3513;
aud[49653]=16'h3507;
aud[49654]=16'h34fb;
aud[49655]=16'h34ef;
aud[49656]=16'h34e3;
aud[49657]=16'h34d7;
aud[49658]=16'h34cb;
aud[49659]=16'h34be;
aud[49660]=16'h34b2;
aud[49661]=16'h34a6;
aud[49662]=16'h349a;
aud[49663]=16'h348e;
aud[49664]=16'h3481;
aud[49665]=16'h3475;
aud[49666]=16'h3469;
aud[49667]=16'h345d;
aud[49668]=16'h3450;
aud[49669]=16'h3444;
aud[49670]=16'h3437;
aud[49671]=16'h342b;
aud[49672]=16'h341f;
aud[49673]=16'h3412;
aud[49674]=16'h3406;
aud[49675]=16'h33f9;
aud[49676]=16'h33ed;
aud[49677]=16'h33e0;
aud[49678]=16'h33d4;
aud[49679]=16'h33c7;
aud[49680]=16'h33ba;
aud[49681]=16'h33ae;
aud[49682]=16'h33a1;
aud[49683]=16'h3394;
aud[49684]=16'h3388;
aud[49685]=16'h337b;
aud[49686]=16'h336e;
aud[49687]=16'h3361;
aud[49688]=16'h3355;
aud[49689]=16'h3348;
aud[49690]=16'h333b;
aud[49691]=16'h332e;
aud[49692]=16'h3321;
aud[49693]=16'h3314;
aud[49694]=16'h3307;
aud[49695]=16'h32fa;
aud[49696]=16'h32ed;
aud[49697]=16'h32e0;
aud[49698]=16'h32d3;
aud[49699]=16'h32c6;
aud[49700]=16'h32b9;
aud[49701]=16'h32ac;
aud[49702]=16'h329f;
aud[49703]=16'h3292;
aud[49704]=16'h3285;
aud[49705]=16'h3278;
aud[49706]=16'h326a;
aud[49707]=16'h325d;
aud[49708]=16'h3250;
aud[49709]=16'h3243;
aud[49710]=16'h3235;
aud[49711]=16'h3228;
aud[49712]=16'h321b;
aud[49713]=16'h320d;
aud[49714]=16'h3200;
aud[49715]=16'h31f3;
aud[49716]=16'h31e5;
aud[49717]=16'h31d8;
aud[49718]=16'h31ca;
aud[49719]=16'h31bd;
aud[49720]=16'h31af;
aud[49721]=16'h31a2;
aud[49722]=16'h3194;
aud[49723]=16'h3187;
aud[49724]=16'h3179;
aud[49725]=16'h316b;
aud[49726]=16'h315e;
aud[49727]=16'h3150;
aud[49728]=16'h3142;
aud[49729]=16'h3135;
aud[49730]=16'h3127;
aud[49731]=16'h3119;
aud[49732]=16'h310b;
aud[49733]=16'h30fe;
aud[49734]=16'h30f0;
aud[49735]=16'h30e2;
aud[49736]=16'h30d4;
aud[49737]=16'h30c6;
aud[49738]=16'h30b8;
aud[49739]=16'h30aa;
aud[49740]=16'h309d;
aud[49741]=16'h308f;
aud[49742]=16'h3081;
aud[49743]=16'h3073;
aud[49744]=16'h3065;
aud[49745]=16'h3057;
aud[49746]=16'h3048;
aud[49747]=16'h303a;
aud[49748]=16'h302c;
aud[49749]=16'h301e;
aud[49750]=16'h3010;
aud[49751]=16'h3002;
aud[49752]=16'h2ff4;
aud[49753]=16'h2fe5;
aud[49754]=16'h2fd7;
aud[49755]=16'h2fc9;
aud[49756]=16'h2fbb;
aud[49757]=16'h2fac;
aud[49758]=16'h2f9e;
aud[49759]=16'h2f90;
aud[49760]=16'h2f81;
aud[49761]=16'h2f73;
aud[49762]=16'h2f65;
aud[49763]=16'h2f56;
aud[49764]=16'h2f48;
aud[49765]=16'h2f39;
aud[49766]=16'h2f2b;
aud[49767]=16'h2f1c;
aud[49768]=16'h2f0e;
aud[49769]=16'h2eff;
aud[49770]=16'h2ef1;
aud[49771]=16'h2ee2;
aud[49772]=16'h2ed3;
aud[49773]=16'h2ec5;
aud[49774]=16'h2eb6;
aud[49775]=16'h2ea7;
aud[49776]=16'h2e99;
aud[49777]=16'h2e8a;
aud[49778]=16'h2e7b;
aud[49779]=16'h2e6d;
aud[49780]=16'h2e5e;
aud[49781]=16'h2e4f;
aud[49782]=16'h2e40;
aud[49783]=16'h2e31;
aud[49784]=16'h2e22;
aud[49785]=16'h2e14;
aud[49786]=16'h2e05;
aud[49787]=16'h2df6;
aud[49788]=16'h2de7;
aud[49789]=16'h2dd8;
aud[49790]=16'h2dc9;
aud[49791]=16'h2dba;
aud[49792]=16'h2dab;
aud[49793]=16'h2d9c;
aud[49794]=16'h2d8d;
aud[49795]=16'h2d7e;
aud[49796]=16'h2d6f;
aud[49797]=16'h2d60;
aud[49798]=16'h2d50;
aud[49799]=16'h2d41;
aud[49800]=16'h2d32;
aud[49801]=16'h2d23;
aud[49802]=16'h2d14;
aud[49803]=16'h2d04;
aud[49804]=16'h2cf5;
aud[49805]=16'h2ce6;
aud[49806]=16'h2cd7;
aud[49807]=16'h2cc7;
aud[49808]=16'h2cb8;
aud[49809]=16'h2ca9;
aud[49810]=16'h2c99;
aud[49811]=16'h2c8a;
aud[49812]=16'h2c7a;
aud[49813]=16'h2c6b;
aud[49814]=16'h2c5c;
aud[49815]=16'h2c4c;
aud[49816]=16'h2c3d;
aud[49817]=16'h2c2d;
aud[49818]=16'h2c1e;
aud[49819]=16'h2c0e;
aud[49820]=16'h2bfe;
aud[49821]=16'h2bef;
aud[49822]=16'h2bdf;
aud[49823]=16'h2bd0;
aud[49824]=16'h2bc0;
aud[49825]=16'h2bb0;
aud[49826]=16'h2ba1;
aud[49827]=16'h2b91;
aud[49828]=16'h2b81;
aud[49829]=16'h2b71;
aud[49830]=16'h2b62;
aud[49831]=16'h2b52;
aud[49832]=16'h2b42;
aud[49833]=16'h2b32;
aud[49834]=16'h2b22;
aud[49835]=16'h2b13;
aud[49836]=16'h2b03;
aud[49837]=16'h2af3;
aud[49838]=16'h2ae3;
aud[49839]=16'h2ad3;
aud[49840]=16'h2ac3;
aud[49841]=16'h2ab3;
aud[49842]=16'h2aa3;
aud[49843]=16'h2a93;
aud[49844]=16'h2a83;
aud[49845]=16'h2a73;
aud[49846]=16'h2a63;
aud[49847]=16'h2a53;
aud[49848]=16'h2a43;
aud[49849]=16'h2a33;
aud[49850]=16'h2a23;
aud[49851]=16'h2a12;
aud[49852]=16'h2a02;
aud[49853]=16'h29f2;
aud[49854]=16'h29e2;
aud[49855]=16'h29d2;
aud[49856]=16'h29c1;
aud[49857]=16'h29b1;
aud[49858]=16'h29a1;
aud[49859]=16'h2991;
aud[49860]=16'h2980;
aud[49861]=16'h2970;
aud[49862]=16'h2960;
aud[49863]=16'h294f;
aud[49864]=16'h293f;
aud[49865]=16'h292e;
aud[49866]=16'h291e;
aud[49867]=16'h290e;
aud[49868]=16'h28fd;
aud[49869]=16'h28ed;
aud[49870]=16'h28dc;
aud[49871]=16'h28cc;
aud[49872]=16'h28bb;
aud[49873]=16'h28aa;
aud[49874]=16'h289a;
aud[49875]=16'h2889;
aud[49876]=16'h2879;
aud[49877]=16'h2868;
aud[49878]=16'h2857;
aud[49879]=16'h2847;
aud[49880]=16'h2836;
aud[49881]=16'h2825;
aud[49882]=16'h2815;
aud[49883]=16'h2804;
aud[49884]=16'h27f3;
aud[49885]=16'h27e2;
aud[49886]=16'h27d2;
aud[49887]=16'h27c1;
aud[49888]=16'h27b0;
aud[49889]=16'h279f;
aud[49890]=16'h278e;
aud[49891]=16'h277e;
aud[49892]=16'h276d;
aud[49893]=16'h275c;
aud[49894]=16'h274b;
aud[49895]=16'h273a;
aud[49896]=16'h2729;
aud[49897]=16'h2718;
aud[49898]=16'h2707;
aud[49899]=16'h26f6;
aud[49900]=16'h26e5;
aud[49901]=16'h26d4;
aud[49902]=16'h26c3;
aud[49903]=16'h26b2;
aud[49904]=16'h26a1;
aud[49905]=16'h2690;
aud[49906]=16'h267e;
aud[49907]=16'h266d;
aud[49908]=16'h265c;
aud[49909]=16'h264b;
aud[49910]=16'h263a;
aud[49911]=16'h2629;
aud[49912]=16'h2617;
aud[49913]=16'h2606;
aud[49914]=16'h25f5;
aud[49915]=16'h25e4;
aud[49916]=16'h25d2;
aud[49917]=16'h25c1;
aud[49918]=16'h25b0;
aud[49919]=16'h259e;
aud[49920]=16'h258d;
aud[49921]=16'h257c;
aud[49922]=16'h256a;
aud[49923]=16'h2559;
aud[49924]=16'h2547;
aud[49925]=16'h2536;
aud[49926]=16'h2524;
aud[49927]=16'h2513;
aud[49928]=16'h2501;
aud[49929]=16'h24f0;
aud[49930]=16'h24de;
aud[49931]=16'h24cd;
aud[49932]=16'h24bb;
aud[49933]=16'h24aa;
aud[49934]=16'h2498;
aud[49935]=16'h2487;
aud[49936]=16'h2475;
aud[49937]=16'h2463;
aud[49938]=16'h2452;
aud[49939]=16'h2440;
aud[49940]=16'h242e;
aud[49941]=16'h241d;
aud[49942]=16'h240b;
aud[49943]=16'h23f9;
aud[49944]=16'h23e7;
aud[49945]=16'h23d6;
aud[49946]=16'h23c4;
aud[49947]=16'h23b2;
aud[49948]=16'h23a0;
aud[49949]=16'h238e;
aud[49950]=16'h237d;
aud[49951]=16'h236b;
aud[49952]=16'h2359;
aud[49953]=16'h2347;
aud[49954]=16'h2335;
aud[49955]=16'h2323;
aud[49956]=16'h2311;
aud[49957]=16'h22ff;
aud[49958]=16'h22ed;
aud[49959]=16'h22db;
aud[49960]=16'h22c9;
aud[49961]=16'h22b7;
aud[49962]=16'h22a5;
aud[49963]=16'h2293;
aud[49964]=16'h2281;
aud[49965]=16'h226f;
aud[49966]=16'h225d;
aud[49967]=16'h224b;
aud[49968]=16'h2239;
aud[49969]=16'h2227;
aud[49970]=16'h2215;
aud[49971]=16'h2202;
aud[49972]=16'h21f0;
aud[49973]=16'h21de;
aud[49974]=16'h21cc;
aud[49975]=16'h21ba;
aud[49976]=16'h21a7;
aud[49977]=16'h2195;
aud[49978]=16'h2183;
aud[49979]=16'h2171;
aud[49980]=16'h215e;
aud[49981]=16'h214c;
aud[49982]=16'h213a;
aud[49983]=16'h2127;
aud[49984]=16'h2115;
aud[49985]=16'h2103;
aud[49986]=16'h20f0;
aud[49987]=16'h20de;
aud[49988]=16'h20cb;
aud[49989]=16'h20b9;
aud[49990]=16'h20a7;
aud[49991]=16'h2094;
aud[49992]=16'h2082;
aud[49993]=16'h206f;
aud[49994]=16'h205d;
aud[49995]=16'h204a;
aud[49996]=16'h2038;
aud[49997]=16'h2025;
aud[49998]=16'h2013;
aud[49999]=16'h2000;

end


endmodule