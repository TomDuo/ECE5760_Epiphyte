module testVect (
output reg signed [15:0] aud [0:1999]
);

initial begin
aud[0]=16'h78;
aud[1]=16'hef;
aud[2]=16'h161;
aud[3]=16'h1cd;
aud[4]=16'h231;
aud[5]=16'h28c;
aud[6]=16'h2db;
aud[7]=16'h31e;
aud[8]=16'h353;
aud[9]=16'h37a;
aud[10]=16'h392;
aud[11]=16'h39a;
aud[12]=16'h392;
aud[13]=16'h37a;
aud[14]=16'h353;
aud[15]=16'h31e;
aud[16]=16'h2db;
aud[17]=16'h28c;
aud[18]=16'h231;
aud[19]=16'h1cd;
aud[20]=16'h161;
aud[21]=16'hef;
aud[22]=16'h78;
aud[23]=16'h0;
aud[24]=16'hff88;
aud[25]=16'hff11;
aud[26]=16'hfe9f;
aud[27]=16'hfe33;
aud[28]=16'hfdcf;
aud[29]=16'hfd74;
aud[30]=16'hfd25;
aud[31]=16'hfce2;
aud[32]=16'hfcad;
aud[33]=16'hfc86;
aud[34]=16'hfc6e;
aud[35]=16'hfc66;
aud[36]=16'hfc6e;
aud[37]=16'hfc86;
aud[38]=16'hfcad;
aud[39]=16'hfce2;
aud[40]=16'hfd25;
aud[41]=16'hfd74;
aud[42]=16'hfdcf;
aud[43]=16'hfe33;
aud[44]=16'hfe9f;
aud[45]=16'hff11;
aud[46]=16'hff88;
aud[47]=16'h0;
aud[48]=16'h78;
aud[49]=16'hef;
aud[50]=16'h161;
aud[51]=16'h1cd;
aud[52]=16'h231;
aud[53]=16'h28c;
aud[54]=16'h2db;
aud[55]=16'h31e;
aud[56]=16'h353;
aud[57]=16'h37a;
aud[58]=16'h392;
aud[59]=16'h39a;
aud[60]=16'h392;
aud[61]=16'h37a;
aud[62]=16'h353;
aud[63]=16'h31e;
aud[64]=16'h2db;
aud[65]=16'h28c;
aud[66]=16'h231;
aud[67]=16'h1cd;
aud[68]=16'h161;
aud[69]=16'hef;
aud[70]=16'h78;
aud[71]=16'h0;
aud[72]=16'hff88;
aud[73]=16'hff11;
aud[74]=16'hfe9f;
aud[75]=16'hfe33;
aud[76]=16'hfdcf;
aud[77]=16'hfd74;
aud[78]=16'hfd25;
aud[79]=16'hfce2;
aud[80]=16'hfcad;
aud[81]=16'hfc86;
aud[82]=16'hfc6e;
aud[83]=16'hfc66;
aud[84]=16'hfc6e;
aud[85]=16'hfc86;
aud[86]=16'hfcad;
aud[87]=16'hfce2;
aud[88]=16'hfd25;
aud[89]=16'hfd74;
aud[90]=16'hfdcf;
aud[91]=16'hfe33;
aud[92]=16'hfe9f;
aud[93]=16'hff11;
aud[94]=16'hff88;
aud[95]=16'h0;
aud[96]=16'h78;
aud[97]=16'hef;
aud[98]=16'h161;
aud[99]=16'h1cd;
aud[100]=16'h231;
aud[101]=16'h28c;
aud[102]=16'h2db;
aud[103]=16'h31e;
aud[104]=16'h353;
aud[105]=16'h37a;
aud[106]=16'h392;
aud[107]=16'h39a;
aud[108]=16'h392;
aud[109]=16'h37a;
aud[110]=16'h353;
aud[111]=16'h31e;
aud[112]=16'h2db;
aud[113]=16'h28c;
aud[114]=16'h231;
aud[115]=16'h1cd;
aud[116]=16'h161;
aud[117]=16'hef;
aud[118]=16'h78;
aud[119]=16'h0;
aud[120]=16'hff88;
aud[121]=16'hff11;
aud[122]=16'hfe9f;
aud[123]=16'hfe33;
aud[124]=16'hfdcf;
aud[125]=16'hfd74;
aud[126]=16'hfd25;
aud[127]=16'hfce2;
aud[128]=16'hfcad;
aud[129]=16'hfc86;
aud[130]=16'hfc6e;
aud[131]=16'hfc66;
aud[132]=16'hfc6e;
aud[133]=16'hfc86;
aud[134]=16'hfcad;
aud[135]=16'hfce2;
aud[136]=16'hfd25;
aud[137]=16'hfd74;
aud[138]=16'hfdcf;
aud[139]=16'hfe33;
aud[140]=16'hfe9f;
aud[141]=16'hff11;
aud[142]=16'hff88;
aud[143]=16'h0;
aud[144]=16'h78;
aud[145]=16'hef;
aud[146]=16'h161;
aud[147]=16'h1cd;
aud[148]=16'h231;
aud[149]=16'h28c;
aud[150]=16'h2db;
aud[151]=16'h31e;
aud[152]=16'h353;
aud[153]=16'h37a;
aud[154]=16'h392;
aud[155]=16'h39a;
aud[156]=16'h392;
aud[157]=16'h37a;
aud[158]=16'h353;
aud[159]=16'h31e;
aud[160]=16'h2db;
aud[161]=16'h28c;
aud[162]=16'h231;
aud[163]=16'h1cd;
aud[164]=16'h161;
aud[165]=16'hef;
aud[166]=16'h78;
aud[167]=16'h0;
aud[168]=16'hff88;
aud[169]=16'hff11;
aud[170]=16'hfe9f;
aud[171]=16'hfe33;
aud[172]=16'hfdcf;
aud[173]=16'hfd74;
aud[174]=16'hfd25;
aud[175]=16'hfce2;
aud[176]=16'hfcad;
aud[177]=16'hfc86;
aud[178]=16'hfc6e;
aud[179]=16'hfc66;
aud[180]=16'hfc6e;
aud[181]=16'hfc86;
aud[182]=16'hfcad;
aud[183]=16'hfce2;
aud[184]=16'hfd25;
aud[185]=16'hfd74;
aud[186]=16'hfdcf;
aud[187]=16'hfe33;
aud[188]=16'hfe9f;
aud[189]=16'hff11;
aud[190]=16'hff88;
aud[191]=16'h0;
aud[192]=16'h78;
aud[193]=16'hef;
aud[194]=16'h161;
aud[195]=16'h1cd;
aud[196]=16'h231;
aud[197]=16'h28c;
aud[198]=16'h2db;
aud[199]=16'h31e;
aud[200]=16'h353;
aud[201]=16'h37a;
aud[202]=16'h392;
aud[203]=16'h39a;
aud[204]=16'h392;
aud[205]=16'h37a;
aud[206]=16'h353;
aud[207]=16'h31e;
aud[208]=16'h2db;
aud[209]=16'h28c;
aud[210]=16'h231;
aud[211]=16'h1cd;
aud[212]=16'h161;
aud[213]=16'hef;
aud[214]=16'h78;
aud[215]=16'h0;
aud[216]=16'hff88;
aud[217]=16'hff11;
aud[218]=16'hfe9f;
aud[219]=16'hfe33;
aud[220]=16'hfdcf;
aud[221]=16'hfd74;
aud[222]=16'hfd25;
aud[223]=16'hfce2;
aud[224]=16'hfcad;
aud[225]=16'hfc86;
aud[226]=16'hfc6e;
aud[227]=16'hfc66;
aud[228]=16'hfc6e;
aud[229]=16'hfc86;
aud[230]=16'hfcad;
aud[231]=16'hfce2;
aud[232]=16'hfd25;
aud[233]=16'hfd74;
aud[234]=16'hfdcf;
aud[235]=16'hfe33;
aud[236]=16'hfe9f;
aud[237]=16'hff11;
aud[238]=16'hff88;
aud[239]=16'h0;
aud[240]=16'h78;
aud[241]=16'hef;
aud[242]=16'h161;
aud[243]=16'h1cd;
aud[244]=16'h231;
aud[245]=16'h28c;
aud[246]=16'h2db;
aud[247]=16'h31e;
aud[248]=16'h353;
aud[249]=16'h37a;
aud[250]=16'h392;
aud[251]=16'h39a;
aud[252]=16'h392;
aud[253]=16'h37a;
aud[254]=16'h353;
aud[255]=16'h31e;
aud[256]=16'h2db;
aud[257]=16'h28c;
aud[258]=16'h231;
aud[259]=16'h1cd;
aud[260]=16'h161;
aud[261]=16'hef;
aud[262]=16'h78;
aud[263]=16'h0;
aud[264]=16'hff88;
aud[265]=16'hff11;
aud[266]=16'hfe9f;
aud[267]=16'hfe33;
aud[268]=16'hfdcf;
aud[269]=16'hfd74;
aud[270]=16'hfd25;
aud[271]=16'hfce2;
aud[272]=16'hfcad;
aud[273]=16'hfc86;
aud[274]=16'hfc6e;
aud[275]=16'hfc66;
aud[276]=16'hfc6e;
aud[277]=16'hfc86;
aud[278]=16'hfcad;
aud[279]=16'hfce2;
aud[280]=16'hfd25;
aud[281]=16'hfd74;
aud[282]=16'hfdcf;
aud[283]=16'hfe33;
aud[284]=16'hfe9f;
aud[285]=16'hff11;
aud[286]=16'hff88;
aud[287]=16'h0;
aud[288]=16'h78;
aud[289]=16'hef;
aud[290]=16'h161;
aud[291]=16'h1cd;
aud[292]=16'h231;
aud[293]=16'h28c;
aud[294]=16'h2db;
aud[295]=16'h31e;
aud[296]=16'h353;
aud[297]=16'h37a;
aud[298]=16'h392;
aud[299]=16'h39a;
aud[300]=16'h392;
aud[301]=16'h37a;
aud[302]=16'h353;
aud[303]=16'h31e;
aud[304]=16'h2db;
aud[305]=16'h28c;
aud[306]=16'h231;
aud[307]=16'h1cd;
aud[308]=16'h161;
aud[309]=16'hef;
aud[310]=16'h78;
aud[311]=16'h0;
aud[312]=16'hff88;
aud[313]=16'hff11;
aud[314]=16'hfe9f;
aud[315]=16'hfe33;
aud[316]=16'hfdcf;
aud[317]=16'hfd74;
aud[318]=16'hfd25;
aud[319]=16'hfce2;
aud[320]=16'hfcad;
aud[321]=16'hfc86;
aud[322]=16'hfc6e;
aud[323]=16'hfc66;
aud[324]=16'hfc6e;
aud[325]=16'hfc86;
aud[326]=16'hfcad;
aud[327]=16'hfce2;
aud[328]=16'hfd25;
aud[329]=16'hfd74;
aud[330]=16'hfdcf;
aud[331]=16'hfe33;
aud[332]=16'hfe9f;
aud[333]=16'hff11;
aud[334]=16'hff88;
aud[335]=16'h0;
aud[336]=16'h78;
aud[337]=16'hef;
aud[338]=16'h161;
aud[339]=16'h1cd;
aud[340]=16'h231;
aud[341]=16'h28c;
aud[342]=16'h2db;
aud[343]=16'h31e;
aud[344]=16'h353;
aud[345]=16'h37a;
aud[346]=16'h392;
aud[347]=16'h39a;
aud[348]=16'h392;
aud[349]=16'h37a;
aud[350]=16'h353;
aud[351]=16'h31e;
aud[352]=16'h2db;
aud[353]=16'h28c;
aud[354]=16'h231;
aud[355]=16'h1cd;
aud[356]=16'h161;
aud[357]=16'hef;
aud[358]=16'h78;
aud[359]=16'h0;
aud[360]=16'hff88;
aud[361]=16'hff11;
aud[362]=16'hfe9f;
aud[363]=16'hfe33;
aud[364]=16'hfdcf;
aud[365]=16'hfd74;
aud[366]=16'hfd25;
aud[367]=16'hfce2;
aud[368]=16'hfcad;
aud[369]=16'hfc86;
aud[370]=16'hfc6e;
aud[371]=16'hfc66;
aud[372]=16'hfc6e;
aud[373]=16'hfc86;
aud[374]=16'hfcad;
aud[375]=16'hfce2;
aud[376]=16'hfd25;
aud[377]=16'hfd74;
aud[378]=16'hfdcf;
aud[379]=16'hfe33;
aud[380]=16'hfe9f;
aud[381]=16'hff11;
aud[382]=16'hff88;
aud[383]=16'h0;
aud[384]=16'h78;
aud[385]=16'hef;
aud[386]=16'h161;
aud[387]=16'h1cd;
aud[388]=16'h231;
aud[389]=16'h28c;
aud[390]=16'h2db;
aud[391]=16'h31e;
aud[392]=16'h353;
aud[393]=16'h37a;
aud[394]=16'h392;
aud[395]=16'h39a;
aud[396]=16'h392;
aud[397]=16'h37a;
aud[398]=16'h353;
aud[399]=16'h31e;
aud[400]=16'h2db;
aud[401]=16'h28c;
aud[402]=16'h231;
aud[403]=16'h1cd;
aud[404]=16'h161;
aud[405]=16'hef;
aud[406]=16'h78;
aud[407]=16'h0;
aud[408]=16'hff88;
aud[409]=16'hff11;
aud[410]=16'hfe9f;
aud[411]=16'hfe33;
aud[412]=16'hfdcf;
aud[413]=16'hfd74;
aud[414]=16'hfd25;
aud[415]=16'hfce2;
aud[416]=16'hfcad;
aud[417]=16'hfc86;
aud[418]=16'hfc6e;
aud[419]=16'hfc66;
aud[420]=16'hfc6e;
aud[421]=16'hfc86;
aud[422]=16'hfcad;
aud[423]=16'hfce2;
aud[424]=16'hfd25;
aud[425]=16'hfd74;
aud[426]=16'hfdcf;
aud[427]=16'hfe33;
aud[428]=16'hfe9f;
aud[429]=16'hff11;
aud[430]=16'hff88;
aud[431]=16'h0;
aud[432]=16'h78;
aud[433]=16'hef;
aud[434]=16'h161;
aud[435]=16'h1cd;
aud[436]=16'h231;
aud[437]=16'h28c;
aud[438]=16'h2db;
aud[439]=16'h31e;
aud[440]=16'h353;
aud[441]=16'h37a;
aud[442]=16'h392;
aud[443]=16'h39a;
aud[444]=16'h392;
aud[445]=16'h37a;
aud[446]=16'h353;
aud[447]=16'h31e;
aud[448]=16'h2db;
aud[449]=16'h28c;
aud[450]=16'h231;
aud[451]=16'h1cd;
aud[452]=16'h161;
aud[453]=16'hef;
aud[454]=16'h78;
aud[455]=16'h0;
aud[456]=16'hff88;
aud[457]=16'hff11;
aud[458]=16'hfe9f;
aud[459]=16'hfe33;
aud[460]=16'hfdcf;
aud[461]=16'hfd74;
aud[462]=16'hfd25;
aud[463]=16'hfce2;
aud[464]=16'hfcad;
aud[465]=16'hfc86;
aud[466]=16'hfc6e;
aud[467]=16'hfc66;
aud[468]=16'hfc6e;
aud[469]=16'hfc86;
aud[470]=16'hfcad;
aud[471]=16'hfce2;
aud[472]=16'hfd25;
aud[473]=16'hfd74;
aud[474]=16'hfdcf;
aud[475]=16'hfe33;
aud[476]=16'hfe9f;
aud[477]=16'hff11;
aud[478]=16'hff88;
aud[479]=16'h0;
aud[480]=16'h78;
aud[481]=16'hef;
aud[482]=16'h161;
aud[483]=16'h1cd;
aud[484]=16'h231;
aud[485]=16'h28c;
aud[486]=16'h2db;
aud[487]=16'h31e;
aud[488]=16'h353;
aud[489]=16'h37a;
aud[490]=16'h392;
aud[491]=16'h39a;
aud[492]=16'h392;
aud[493]=16'h37a;
aud[494]=16'h353;
aud[495]=16'h31e;
aud[496]=16'h2db;
aud[497]=16'h28c;
aud[498]=16'h231;
aud[499]=16'h1cd;
aud[500]=16'h161;
aud[501]=16'hef;
aud[502]=16'h78;
aud[503]=16'h0;
aud[504]=16'hff88;
aud[505]=16'hff11;
aud[506]=16'hfe9f;
aud[507]=16'hfe33;
aud[508]=16'hfdcf;
aud[509]=16'hfd74;
aud[510]=16'hfd25;
aud[511]=16'hfce2;
aud[512]=16'hfcad;
aud[513]=16'hfc86;
aud[514]=16'hfc6e;
aud[515]=16'hfc66;
aud[516]=16'hfc6e;
aud[517]=16'hfc86;
aud[518]=16'hfcad;
aud[519]=16'hfce2;
aud[520]=16'hfd25;
aud[521]=16'hfd74;
aud[522]=16'hfdcf;
aud[523]=16'hfe33;
aud[524]=16'hfe9f;
aud[525]=16'hff11;
aud[526]=16'hff88;
aud[527]=16'h0;
aud[528]=16'h78;
aud[529]=16'hef;
aud[530]=16'h161;
aud[531]=16'h1cd;
aud[532]=16'h231;
aud[533]=16'h28c;
aud[534]=16'h2db;
aud[535]=16'h31e;
aud[536]=16'h353;
aud[537]=16'h37a;
aud[538]=16'h392;
aud[539]=16'h39a;
aud[540]=16'h392;
aud[541]=16'h37a;
aud[542]=16'h353;
aud[543]=16'h31e;
aud[544]=16'h2db;
aud[545]=16'h28c;
aud[546]=16'h231;
aud[547]=16'h1cd;
aud[548]=16'h161;
aud[549]=16'hef;
aud[550]=16'h78;
aud[551]=16'h0;
aud[552]=16'hff88;
aud[553]=16'hff11;
aud[554]=16'hfe9f;
aud[555]=16'hfe33;
aud[556]=16'hfdcf;
aud[557]=16'hfd74;
aud[558]=16'hfd25;
aud[559]=16'hfce2;
aud[560]=16'hfcad;
aud[561]=16'hfc86;
aud[562]=16'hfc6e;
aud[563]=16'hfc66;
aud[564]=16'hfc6e;
aud[565]=16'hfc86;
aud[566]=16'hfcad;
aud[567]=16'hfce2;
aud[568]=16'hfd25;
aud[569]=16'hfd74;
aud[570]=16'hfdcf;
aud[571]=16'hfe33;
aud[572]=16'hfe9f;
aud[573]=16'hff11;
aud[574]=16'hff88;
aud[575]=16'h0;
aud[576]=16'h78;
aud[577]=16'hef;
aud[578]=16'h161;
aud[579]=16'h1cd;
aud[580]=16'h231;
aud[581]=16'h28c;
aud[582]=16'h2db;
aud[583]=16'h31e;
aud[584]=16'h353;
aud[585]=16'h37a;
aud[586]=16'h392;
aud[587]=16'h39a;
aud[588]=16'h392;
aud[589]=16'h37a;
aud[590]=16'h353;
aud[591]=16'h31e;
aud[592]=16'h2db;
aud[593]=16'h28c;
aud[594]=16'h231;
aud[595]=16'h1cd;
aud[596]=16'h161;
aud[597]=16'hef;
aud[598]=16'h78;
aud[599]=16'h0;
aud[600]=16'hff88;
aud[601]=16'hff11;
aud[602]=16'hfe9f;
aud[603]=16'hfe33;
aud[604]=16'hfdcf;
aud[605]=16'hfd74;
aud[606]=16'hfd25;
aud[607]=16'hfce2;
aud[608]=16'hfcad;
aud[609]=16'hfc86;
aud[610]=16'hfc6e;
aud[611]=16'hfc66;
aud[612]=16'hfc6e;
aud[613]=16'hfc86;
aud[614]=16'hfcad;
aud[615]=16'hfce2;
aud[616]=16'hfd25;
aud[617]=16'hfd74;
aud[618]=16'hfdcf;
aud[619]=16'hfe33;
aud[620]=16'hfe9f;
aud[621]=16'hff11;
aud[622]=16'hff88;
aud[623]=16'h0;
aud[624]=16'h78;
aud[625]=16'hef;
aud[626]=16'h161;
aud[627]=16'h1cd;
aud[628]=16'h231;
aud[629]=16'h28c;
aud[630]=16'h2db;
aud[631]=16'h31e;
aud[632]=16'h353;
aud[633]=16'h37a;
aud[634]=16'h392;
aud[635]=16'h39a;
aud[636]=16'h392;
aud[637]=16'h37a;
aud[638]=16'h353;
aud[639]=16'h31e;
aud[640]=16'h2db;
aud[641]=16'h28c;
aud[642]=16'h231;
aud[643]=16'h1cd;
aud[644]=16'h161;
aud[645]=16'hef;
aud[646]=16'h78;
aud[647]=16'h0;
aud[648]=16'hff88;
aud[649]=16'hff11;
aud[650]=16'hfe9f;
aud[651]=16'hfe33;
aud[652]=16'hfdcf;
aud[653]=16'hfd74;
aud[654]=16'hfd25;
aud[655]=16'hfce2;
aud[656]=16'hfcad;
aud[657]=16'hfc86;
aud[658]=16'hfc6e;
aud[659]=16'hfc66;
aud[660]=16'hfc6e;
aud[661]=16'hfc86;
aud[662]=16'hfcad;
aud[663]=16'hfce2;
aud[664]=16'hfd25;
aud[665]=16'hfd74;
aud[666]=16'hfdcf;
aud[667]=16'hfe33;
aud[668]=16'hfe9f;
aud[669]=16'hff11;
aud[670]=16'hff88;
aud[671]=16'h0;
aud[672]=16'h78;
aud[673]=16'hef;
aud[674]=16'h161;
aud[675]=16'h1cd;
aud[676]=16'h231;
aud[677]=16'h28c;
aud[678]=16'h2db;
aud[679]=16'h31e;
aud[680]=16'h353;
aud[681]=16'h37a;
aud[682]=16'h392;
aud[683]=16'h39a;
aud[684]=16'h392;
aud[685]=16'h37a;
aud[686]=16'h353;
aud[687]=16'h31e;
aud[688]=16'h2db;
aud[689]=16'h28c;
aud[690]=16'h231;
aud[691]=16'h1cd;
aud[692]=16'h161;
aud[693]=16'hef;
aud[694]=16'h78;
aud[695]=16'h0;
aud[696]=16'hff88;
aud[697]=16'hff11;
aud[698]=16'hfe9f;
aud[699]=16'hfe33;
aud[700]=16'hfdcf;
aud[701]=16'hfd74;
aud[702]=16'hfd25;
aud[703]=16'hfce2;
aud[704]=16'hfcad;
aud[705]=16'hfc86;
aud[706]=16'hfc6e;
aud[707]=16'hfc66;
aud[708]=16'hfc6e;
aud[709]=16'hfc86;
aud[710]=16'hfcad;
aud[711]=16'hfce2;
aud[712]=16'hfd25;
aud[713]=16'hfd74;
aud[714]=16'hfdcf;
aud[715]=16'hfe33;
aud[716]=16'hfe9f;
aud[717]=16'hff11;
aud[718]=16'hff88;
aud[719]=16'h0;
aud[720]=16'h78;
aud[721]=16'hef;
aud[722]=16'h161;
aud[723]=16'h1cd;
aud[724]=16'h231;
aud[725]=16'h28c;
aud[726]=16'h2db;
aud[727]=16'h31e;
aud[728]=16'h353;
aud[729]=16'h37a;
aud[730]=16'h392;
aud[731]=16'h39a;
aud[732]=16'h392;
aud[733]=16'h37a;
aud[734]=16'h353;
aud[735]=16'h31e;
aud[736]=16'h2db;
aud[737]=16'h28c;
aud[738]=16'h231;
aud[739]=16'h1cd;
aud[740]=16'h161;
aud[741]=16'hef;
aud[742]=16'h78;
aud[743]=16'h0;
aud[744]=16'hff88;
aud[745]=16'hff11;
aud[746]=16'hfe9f;
aud[747]=16'hfe33;
aud[748]=16'hfdcf;
aud[749]=16'hfd74;
aud[750]=16'hfd25;
aud[751]=16'hfce2;
aud[752]=16'hfcad;
aud[753]=16'hfc86;
aud[754]=16'hfc6e;
aud[755]=16'hfc66;
aud[756]=16'hfc6e;
aud[757]=16'hfc86;
aud[758]=16'hfcad;
aud[759]=16'hfce2;
aud[760]=16'hfd25;
aud[761]=16'hfd74;
aud[762]=16'hfdcf;
aud[763]=16'hfe33;
aud[764]=16'hfe9f;
aud[765]=16'hff11;
aud[766]=16'hff88;
aud[767]=16'h0;
aud[768]=16'h78;
aud[769]=16'hef;
aud[770]=16'h161;
aud[771]=16'h1cd;
aud[772]=16'h231;
aud[773]=16'h28c;
aud[774]=16'h2db;
aud[775]=16'h31e;
aud[776]=16'h353;
aud[777]=16'h37a;
aud[778]=16'h392;
aud[779]=16'h39a;
aud[780]=16'h392;
aud[781]=16'h37a;
aud[782]=16'h353;
aud[783]=16'h31e;
aud[784]=16'h2db;
aud[785]=16'h28c;
aud[786]=16'h231;
aud[787]=16'h1cd;
aud[788]=16'h161;
aud[789]=16'hef;
aud[790]=16'h78;
aud[791]=16'h0;
aud[792]=16'hff88;
aud[793]=16'hff11;
aud[794]=16'hfe9f;
aud[795]=16'hfe33;
aud[796]=16'hfdcf;
aud[797]=16'hfd74;
aud[798]=16'hfd25;
aud[799]=16'hfce2;
aud[800]=16'hfcad;
aud[801]=16'hfc86;
aud[802]=16'hfc6e;
aud[803]=16'hfc66;
aud[804]=16'hfc6e;
aud[805]=16'hfc86;
aud[806]=16'hfcad;
aud[807]=16'hfce2;
aud[808]=16'hfd25;
aud[809]=16'hfd74;
aud[810]=16'hfdcf;
aud[811]=16'hfe33;
aud[812]=16'hfe9f;
aud[813]=16'hff11;
aud[814]=16'hff88;
aud[815]=16'h0;
aud[816]=16'h78;
aud[817]=16'hef;
aud[818]=16'h161;
aud[819]=16'h1cd;
aud[820]=16'h231;
aud[821]=16'h28c;
aud[822]=16'h2db;
aud[823]=16'h31e;
aud[824]=16'h353;
aud[825]=16'h37a;
aud[826]=16'h392;
aud[827]=16'h39a;
aud[828]=16'h392;
aud[829]=16'h37a;
aud[830]=16'h353;
aud[831]=16'h31e;
aud[832]=16'h2db;
aud[833]=16'h28c;
aud[834]=16'h231;
aud[835]=16'h1cd;
aud[836]=16'h161;
aud[837]=16'hef;
aud[838]=16'h78;
aud[839]=16'h0;
aud[840]=16'hff88;
aud[841]=16'hff11;
aud[842]=16'hfe9f;
aud[843]=16'hfe33;
aud[844]=16'hfdcf;
aud[845]=16'hfd74;
aud[846]=16'hfd25;
aud[847]=16'hfce2;
aud[848]=16'hfcad;
aud[849]=16'hfc86;
aud[850]=16'hfc6e;
aud[851]=16'hfc66;
aud[852]=16'hfc6e;
aud[853]=16'hfc86;
aud[854]=16'hfcad;
aud[855]=16'hfce2;
aud[856]=16'hfd25;
aud[857]=16'hfd74;
aud[858]=16'hfdcf;
aud[859]=16'hfe33;
aud[860]=16'hfe9f;
aud[861]=16'hff11;
aud[862]=16'hff88;
aud[863]=16'h0;
aud[864]=16'h78;
aud[865]=16'hef;
aud[866]=16'h161;
aud[867]=16'h1cd;
aud[868]=16'h231;
aud[869]=16'h28c;
aud[870]=16'h2db;
aud[871]=16'h31e;
aud[872]=16'h353;
aud[873]=16'h37a;
aud[874]=16'h392;
aud[875]=16'h39a;
aud[876]=16'h392;
aud[877]=16'h37a;
aud[878]=16'h353;
aud[879]=16'h31e;
aud[880]=16'h2db;
aud[881]=16'h28c;
aud[882]=16'h231;
aud[883]=16'h1cd;
aud[884]=16'h161;
aud[885]=16'hef;
aud[886]=16'h78;
aud[887]=16'h0;
aud[888]=16'hff88;
aud[889]=16'hff11;
aud[890]=16'hfe9f;
aud[891]=16'hfe33;
aud[892]=16'hfdcf;
aud[893]=16'hfd74;
aud[894]=16'hfd25;
aud[895]=16'hfce2;
aud[896]=16'hfcad;
aud[897]=16'hfc86;
aud[898]=16'hfc6e;
aud[899]=16'hfc66;
aud[900]=16'hfc6e;
aud[901]=16'hfc86;
aud[902]=16'hfcad;
aud[903]=16'hfce2;
aud[904]=16'hfd25;
aud[905]=16'hfd74;
aud[906]=16'hfdcf;
aud[907]=16'hfe33;
aud[908]=16'hfe9f;
aud[909]=16'hff11;
aud[910]=16'hff88;
aud[911]=16'h0;
aud[912]=16'h78;
aud[913]=16'hef;
aud[914]=16'h161;
aud[915]=16'h1cd;
aud[916]=16'h231;
aud[917]=16'h28c;
aud[918]=16'h2db;
aud[919]=16'h31e;
aud[920]=16'h353;
aud[921]=16'h37a;
aud[922]=16'h392;
aud[923]=16'h39a;
aud[924]=16'h392;
aud[925]=16'h37a;
aud[926]=16'h353;
aud[927]=16'h31e;
aud[928]=16'h2db;
aud[929]=16'h28c;
aud[930]=16'h231;
aud[931]=16'h1cd;
aud[932]=16'h161;
aud[933]=16'hef;
aud[934]=16'h78;
aud[935]=16'h0;
aud[936]=16'hff88;
aud[937]=16'hff11;
aud[938]=16'hfe9f;
aud[939]=16'hfe33;
aud[940]=16'hfdcf;
aud[941]=16'hfd74;
aud[942]=16'hfd25;
aud[943]=16'hfce2;
aud[944]=16'hfcad;
aud[945]=16'hfc86;
aud[946]=16'hfc6e;
aud[947]=16'hfc66;
aud[948]=16'hfc6e;
aud[949]=16'hfc86;
aud[950]=16'hfcad;
aud[951]=16'hfce2;
aud[952]=16'hfd25;
aud[953]=16'hfd74;
aud[954]=16'hfdcf;
aud[955]=16'hfe33;
aud[956]=16'hfe9f;
aud[957]=16'hff11;
aud[958]=16'hff88;
aud[959]=16'h0;
aud[960]=16'h78;
aud[961]=16'hef;
aud[962]=16'h161;
aud[963]=16'h1cd;
aud[964]=16'h231;
aud[965]=16'h28c;
aud[966]=16'h2db;
aud[967]=16'h31e;
aud[968]=16'h353;
aud[969]=16'h37a;
aud[970]=16'h392;
aud[971]=16'h39a;
aud[972]=16'h392;
aud[973]=16'h37a;
aud[974]=16'h353;
aud[975]=16'h31e;
aud[976]=16'h2db;
aud[977]=16'h28c;
aud[978]=16'h231;
aud[979]=16'h1cd;
aud[980]=16'h161;
aud[981]=16'hef;
aud[982]=16'h78;
aud[983]=16'h0;
aud[984]=16'hff88;
aud[985]=16'hff11;
aud[986]=16'hfe9f;
aud[987]=16'hfe33;
aud[988]=16'hfdcf;
aud[989]=16'hfd74;
aud[990]=16'hfd25;
aud[991]=16'hfce2;
aud[992]=16'hfcad;
aud[993]=16'hfc86;
aud[994]=16'hfc6e;
aud[995]=16'hfc66;
aud[996]=16'hfc6e;
aud[997]=16'hfc86;
aud[998]=16'hfcad;
aud[999]=16'hfce2;
aud[1000]=16'hfd25;
aud[1001]=16'hfd74;
aud[1002]=16'hfdcf;
aud[1003]=16'hfe33;
aud[1004]=16'hfe9f;
aud[1005]=16'hff11;
aud[1006]=16'hff88;
aud[1007]=16'h0;
aud[1008]=16'h78;
aud[1009]=16'hef;
aud[1010]=16'h161;
aud[1011]=16'h1cd;
aud[1012]=16'h231;
aud[1013]=16'h28c;
aud[1014]=16'h2db;
aud[1015]=16'h31e;
aud[1016]=16'h353;
aud[1017]=16'h37a;
aud[1018]=16'h392;
aud[1019]=16'h39a;
aud[1020]=16'h392;
aud[1021]=16'h37a;
aud[1022]=16'h353;
aud[1023]=16'h31e;
aud[1024]=16'h2db;
aud[1025]=16'h28c;
aud[1026]=16'h231;
aud[1027]=16'h1cd;
aud[1028]=16'h161;
aud[1029]=16'hef;
aud[1030]=16'h78;
aud[1031]=16'h0;
aud[1032]=16'hff88;
aud[1033]=16'hff11;
aud[1034]=16'hfe9f;
aud[1035]=16'hfe33;
aud[1036]=16'hfdcf;
aud[1037]=16'hfd74;
aud[1038]=16'hfd25;
aud[1039]=16'hfce2;
aud[1040]=16'hfcad;
aud[1041]=16'hfc86;
aud[1042]=16'hfc6e;
aud[1043]=16'hfc66;
aud[1044]=16'hfc6e;
aud[1045]=16'hfc86;
aud[1046]=16'hfcad;
aud[1047]=16'hfce2;
aud[1048]=16'hfd25;
aud[1049]=16'hfd74;
aud[1050]=16'hfdcf;
aud[1051]=16'hfe33;
aud[1052]=16'hfe9f;
aud[1053]=16'hff11;
aud[1054]=16'hff88;
aud[1055]=16'h0;
aud[1056]=16'h78;
aud[1057]=16'hef;
aud[1058]=16'h161;
aud[1059]=16'h1cd;
aud[1060]=16'h231;
aud[1061]=16'h28c;
aud[1062]=16'h2db;
aud[1063]=16'h31e;
aud[1064]=16'h353;
aud[1065]=16'h37a;
aud[1066]=16'h392;
aud[1067]=16'h39a;
aud[1068]=16'h392;
aud[1069]=16'h37a;
aud[1070]=16'h353;
aud[1071]=16'h31e;
aud[1072]=16'h2db;
aud[1073]=16'h28c;
aud[1074]=16'h231;
aud[1075]=16'h1cd;
aud[1076]=16'h161;
aud[1077]=16'hef;
aud[1078]=16'h78;
aud[1079]=16'h0;
aud[1080]=16'hff88;
aud[1081]=16'hff11;
aud[1082]=16'hfe9f;
aud[1083]=16'hfe33;
aud[1084]=16'hfdcf;
aud[1085]=16'hfd74;
aud[1086]=16'hfd25;
aud[1087]=16'hfce2;
aud[1088]=16'hfcad;
aud[1089]=16'hfc86;
aud[1090]=16'hfc6e;
aud[1091]=16'hfc66;
aud[1092]=16'hfc6e;
aud[1093]=16'hfc86;
aud[1094]=16'hfcad;
aud[1095]=16'hfce2;
aud[1096]=16'hfd25;
aud[1097]=16'hfd74;
aud[1098]=16'hfdcf;
aud[1099]=16'hfe33;
aud[1100]=16'hfe9f;
aud[1101]=16'hff11;
aud[1102]=16'hff88;
aud[1103]=16'h0;
aud[1104]=16'h78;
aud[1105]=16'hef;
aud[1106]=16'h161;
aud[1107]=16'h1cd;
aud[1108]=16'h231;
aud[1109]=16'h28c;
aud[1110]=16'h2db;
aud[1111]=16'h31e;
aud[1112]=16'h353;
aud[1113]=16'h37a;
aud[1114]=16'h392;
aud[1115]=16'h39a;
aud[1116]=16'h392;
aud[1117]=16'h37a;
aud[1118]=16'h353;
aud[1119]=16'h31e;
aud[1120]=16'h2db;
aud[1121]=16'h28c;
aud[1122]=16'h231;
aud[1123]=16'h1cd;
aud[1124]=16'h161;
aud[1125]=16'hef;
aud[1126]=16'h78;
aud[1127]=16'h0;
aud[1128]=16'hff88;
aud[1129]=16'hff11;
aud[1130]=16'hfe9f;
aud[1131]=16'hfe33;
aud[1132]=16'hfdcf;
aud[1133]=16'hfd74;
aud[1134]=16'hfd25;
aud[1135]=16'hfce2;
aud[1136]=16'hfcad;
aud[1137]=16'hfc86;
aud[1138]=16'hfc6e;
aud[1139]=16'hfc66;
aud[1140]=16'hfc6e;
aud[1141]=16'hfc86;
aud[1142]=16'hfcad;
aud[1143]=16'hfce2;
aud[1144]=16'hfd25;
aud[1145]=16'hfd74;
aud[1146]=16'hfdcf;
aud[1147]=16'hfe33;
aud[1148]=16'hfe9f;
aud[1149]=16'hff11;
aud[1150]=16'hff88;
aud[1151]=16'h0;
aud[1152]=16'h78;
aud[1153]=16'hef;
aud[1154]=16'h161;
aud[1155]=16'h1cd;
aud[1156]=16'h231;
aud[1157]=16'h28c;
aud[1158]=16'h2db;
aud[1159]=16'h31e;
aud[1160]=16'h353;
aud[1161]=16'h37a;
aud[1162]=16'h392;
aud[1163]=16'h39a;
aud[1164]=16'h392;
aud[1165]=16'h37a;
aud[1166]=16'h353;
aud[1167]=16'h31e;
aud[1168]=16'h2db;
aud[1169]=16'h28c;
aud[1170]=16'h231;
aud[1171]=16'h1cd;
aud[1172]=16'h161;
aud[1173]=16'hef;
aud[1174]=16'h78;
aud[1175]=16'h0;
aud[1176]=16'hff88;
aud[1177]=16'hff11;
aud[1178]=16'hfe9f;
aud[1179]=16'hfe33;
aud[1180]=16'hfdcf;
aud[1181]=16'hfd74;
aud[1182]=16'hfd25;
aud[1183]=16'hfce2;
aud[1184]=16'hfcad;
aud[1185]=16'hfc86;
aud[1186]=16'hfc6e;
aud[1187]=16'hfc66;
aud[1188]=16'hfc6e;
aud[1189]=16'hfc86;
aud[1190]=16'hfcad;
aud[1191]=16'hfce2;
aud[1192]=16'hfd25;
aud[1193]=16'hfd74;
aud[1194]=16'hfdcf;
aud[1195]=16'hfe33;
aud[1196]=16'hfe9f;
aud[1197]=16'hff11;
aud[1198]=16'hff88;
aud[1199]=16'h0;
aud[1200]=16'h78;
aud[1201]=16'hef;
aud[1202]=16'h161;
aud[1203]=16'h1cd;
aud[1204]=16'h231;
aud[1205]=16'h28c;
aud[1206]=16'h2db;
aud[1207]=16'h31e;
aud[1208]=16'h353;
aud[1209]=16'h37a;
aud[1210]=16'h392;
aud[1211]=16'h39a;
aud[1212]=16'h392;
aud[1213]=16'h37a;
aud[1214]=16'h353;
aud[1215]=16'h31e;
aud[1216]=16'h2db;
aud[1217]=16'h28c;
aud[1218]=16'h231;
aud[1219]=16'h1cd;
aud[1220]=16'h161;
aud[1221]=16'hef;
aud[1222]=16'h78;
aud[1223]=16'h0;
aud[1224]=16'hff88;
aud[1225]=16'hff11;
aud[1226]=16'hfe9f;
aud[1227]=16'hfe33;
aud[1228]=16'hfdcf;
aud[1229]=16'hfd74;
aud[1230]=16'hfd25;
aud[1231]=16'hfce2;
aud[1232]=16'hfcad;
aud[1233]=16'hfc86;
aud[1234]=16'hfc6e;
aud[1235]=16'hfc66;
aud[1236]=16'hfc6e;
aud[1237]=16'hfc86;
aud[1238]=16'hfcad;
aud[1239]=16'hfce2;
aud[1240]=16'hfd25;
aud[1241]=16'hfd74;
aud[1242]=16'hfdcf;
aud[1243]=16'hfe33;
aud[1244]=16'hfe9f;
aud[1245]=16'hff11;
aud[1246]=16'hff88;
aud[1247]=16'h0;
aud[1248]=16'h78;
aud[1249]=16'hef;
aud[1250]=16'h161;
aud[1251]=16'h1cd;
aud[1252]=16'h231;
aud[1253]=16'h28c;
aud[1254]=16'h2db;
aud[1255]=16'h31e;
aud[1256]=16'h353;
aud[1257]=16'h37a;
aud[1258]=16'h392;
aud[1259]=16'h39a;
aud[1260]=16'h392;
aud[1261]=16'h37a;
aud[1262]=16'h353;
aud[1263]=16'h31e;
aud[1264]=16'h2db;
aud[1265]=16'h28c;
aud[1266]=16'h231;
aud[1267]=16'h1cd;
aud[1268]=16'h161;
aud[1269]=16'hef;
aud[1270]=16'h78;
aud[1271]=16'h0;
aud[1272]=16'hff88;
aud[1273]=16'hff11;
aud[1274]=16'hfe9f;
aud[1275]=16'hfe33;
aud[1276]=16'hfdcf;
aud[1277]=16'hfd74;
aud[1278]=16'hfd25;
aud[1279]=16'hfce2;
aud[1280]=16'hfcad;
aud[1281]=16'hfc86;
aud[1282]=16'hfc6e;
aud[1283]=16'hfc66;
aud[1284]=16'hfc6e;
aud[1285]=16'hfc86;
aud[1286]=16'hfcad;
aud[1287]=16'hfce2;
aud[1288]=16'hfd25;
aud[1289]=16'hfd74;
aud[1290]=16'hfdcf;
aud[1291]=16'hfe33;
aud[1292]=16'hfe9f;
aud[1293]=16'hff11;
aud[1294]=16'hff88;
aud[1295]=16'h0;
aud[1296]=16'h78;
aud[1297]=16'hef;
aud[1298]=16'h161;
aud[1299]=16'h1cd;
aud[1300]=16'h231;
aud[1301]=16'h28c;
aud[1302]=16'h2db;
aud[1303]=16'h31e;
aud[1304]=16'h353;
aud[1305]=16'h37a;
aud[1306]=16'h392;
aud[1307]=16'h39a;
aud[1308]=16'h392;
aud[1309]=16'h37a;
aud[1310]=16'h353;
aud[1311]=16'h31e;
aud[1312]=16'h2db;
aud[1313]=16'h28c;
aud[1314]=16'h231;
aud[1315]=16'h1cd;
aud[1316]=16'h161;
aud[1317]=16'hef;
aud[1318]=16'h78;
aud[1319]=16'h0;
aud[1320]=16'hff88;
aud[1321]=16'hff11;
aud[1322]=16'hfe9f;
aud[1323]=16'hfe33;
aud[1324]=16'hfdcf;
aud[1325]=16'hfd74;
aud[1326]=16'hfd25;
aud[1327]=16'hfce2;
aud[1328]=16'hfcad;
aud[1329]=16'hfc86;
aud[1330]=16'hfc6e;
aud[1331]=16'hfc66;
aud[1332]=16'hfc6e;
aud[1333]=16'hfc86;
aud[1334]=16'hfcad;
aud[1335]=16'hfce2;
aud[1336]=16'hfd25;
aud[1337]=16'hfd74;
aud[1338]=16'hfdcf;
aud[1339]=16'hfe33;
aud[1340]=16'hfe9f;
aud[1341]=16'hff11;
aud[1342]=16'hff88;
aud[1343]=16'h0;
aud[1344]=16'h78;
aud[1345]=16'hef;
aud[1346]=16'h161;
aud[1347]=16'h1cd;
aud[1348]=16'h231;
aud[1349]=16'h28c;
aud[1350]=16'h2db;
aud[1351]=16'h31e;
aud[1352]=16'h353;
aud[1353]=16'h37a;
aud[1354]=16'h392;
aud[1355]=16'h39a;
aud[1356]=16'h392;
aud[1357]=16'h37a;
aud[1358]=16'h353;
aud[1359]=16'h31e;
aud[1360]=16'h2db;
aud[1361]=16'h28c;
aud[1362]=16'h231;
aud[1363]=16'h1cd;
aud[1364]=16'h161;
aud[1365]=16'hef;
aud[1366]=16'h78;
aud[1367]=16'h0;
aud[1368]=16'hff88;
aud[1369]=16'hff11;
aud[1370]=16'hfe9f;
aud[1371]=16'hfe33;
aud[1372]=16'hfdcf;
aud[1373]=16'hfd74;
aud[1374]=16'hfd25;
aud[1375]=16'hfce2;
aud[1376]=16'hfcad;
aud[1377]=16'hfc86;
aud[1378]=16'hfc6e;
aud[1379]=16'hfc66;
aud[1380]=16'hfc6e;
aud[1381]=16'hfc86;
aud[1382]=16'hfcad;
aud[1383]=16'hfce2;
aud[1384]=16'hfd25;
aud[1385]=16'hfd74;
aud[1386]=16'hfdcf;
aud[1387]=16'hfe33;
aud[1388]=16'hfe9f;
aud[1389]=16'hff11;
aud[1390]=16'hff88;
aud[1391]=16'h0;
aud[1392]=16'h78;
aud[1393]=16'hef;
aud[1394]=16'h161;
aud[1395]=16'h1cd;
aud[1396]=16'h231;
aud[1397]=16'h28c;
aud[1398]=16'h2db;
aud[1399]=16'h31e;
aud[1400]=16'h353;
aud[1401]=16'h37a;
aud[1402]=16'h392;
aud[1403]=16'h39a;
aud[1404]=16'h392;
aud[1405]=16'h37a;
aud[1406]=16'h353;
aud[1407]=16'h31e;
aud[1408]=16'h2db;
aud[1409]=16'h28c;
aud[1410]=16'h231;
aud[1411]=16'h1cd;
aud[1412]=16'h161;
aud[1413]=16'hef;
aud[1414]=16'h78;
aud[1415]=16'h0;
aud[1416]=16'hff88;
aud[1417]=16'hff11;
aud[1418]=16'hfe9f;
aud[1419]=16'hfe33;
aud[1420]=16'hfdcf;
aud[1421]=16'hfd74;
aud[1422]=16'hfd25;
aud[1423]=16'hfce2;
aud[1424]=16'hfcad;
aud[1425]=16'hfc86;
aud[1426]=16'hfc6e;
aud[1427]=16'hfc66;
aud[1428]=16'hfc6e;
aud[1429]=16'hfc86;
aud[1430]=16'hfcad;
aud[1431]=16'hfce2;
aud[1432]=16'hfd25;
aud[1433]=16'hfd74;
aud[1434]=16'hfdcf;
aud[1435]=16'hfe33;
aud[1436]=16'hfe9f;
aud[1437]=16'hff11;
aud[1438]=16'hff88;
aud[1439]=16'h0;
aud[1440]=16'h78;
aud[1441]=16'hef;
aud[1442]=16'h161;
aud[1443]=16'h1cd;
aud[1444]=16'h231;
aud[1445]=16'h28c;
aud[1446]=16'h2db;
aud[1447]=16'h31e;
aud[1448]=16'h353;
aud[1449]=16'h37a;
aud[1450]=16'h392;
aud[1451]=16'h39a;
aud[1452]=16'h392;
aud[1453]=16'h37a;
aud[1454]=16'h353;
aud[1455]=16'h31e;
aud[1456]=16'h2db;
aud[1457]=16'h28c;
aud[1458]=16'h231;
aud[1459]=16'h1cd;
aud[1460]=16'h161;
aud[1461]=16'hef;
aud[1462]=16'h78;
aud[1463]=16'h0;
aud[1464]=16'hff88;
aud[1465]=16'hff11;
aud[1466]=16'hfe9f;
aud[1467]=16'hfe33;
aud[1468]=16'hfdcf;
aud[1469]=16'hfd74;
aud[1470]=16'hfd25;
aud[1471]=16'hfce2;
aud[1472]=16'hfcad;
aud[1473]=16'hfc86;
aud[1474]=16'hfc6e;
aud[1475]=16'hfc66;
aud[1476]=16'hfc6e;
aud[1477]=16'hfc86;
aud[1478]=16'hfcad;
aud[1479]=16'hfce2;
aud[1480]=16'hfd25;
aud[1481]=16'hfd74;
aud[1482]=16'hfdcf;
aud[1483]=16'hfe33;
aud[1484]=16'hfe9f;
aud[1485]=16'hff11;
aud[1486]=16'hff88;
aud[1487]=16'h0;
aud[1488]=16'h78;
aud[1489]=16'hef;
aud[1490]=16'h161;
aud[1491]=16'h1cd;
aud[1492]=16'h231;
aud[1493]=16'h28c;
aud[1494]=16'h2db;
aud[1495]=16'h31e;
aud[1496]=16'h353;
aud[1497]=16'h37a;
aud[1498]=16'h392;
aud[1499]=16'h39a;
aud[1500]=16'h392;
aud[1501]=16'h37a;
aud[1502]=16'h353;
aud[1503]=16'h31e;
aud[1504]=16'h2db;
aud[1505]=16'h28c;
aud[1506]=16'h231;
aud[1507]=16'h1cd;
aud[1508]=16'h161;
aud[1509]=16'hef;
aud[1510]=16'h78;
aud[1511]=16'h0;
aud[1512]=16'hff88;
aud[1513]=16'hff11;
aud[1514]=16'hfe9f;
aud[1515]=16'hfe33;
aud[1516]=16'hfdcf;
aud[1517]=16'hfd74;
aud[1518]=16'hfd25;
aud[1519]=16'hfce2;
aud[1520]=16'hfcad;
aud[1521]=16'hfc86;
aud[1522]=16'hfc6e;
aud[1523]=16'hfc66;
aud[1524]=16'hfc6e;
aud[1525]=16'hfc86;
aud[1526]=16'hfcad;
aud[1527]=16'hfce2;
aud[1528]=16'hfd25;
aud[1529]=16'hfd74;
aud[1530]=16'hfdcf;
aud[1531]=16'hfe33;
aud[1532]=16'hfe9f;
aud[1533]=16'hff11;
aud[1534]=16'hff88;
aud[1535]=16'h0;
aud[1536]=16'h78;
aud[1537]=16'hef;
aud[1538]=16'h161;
aud[1539]=16'h1cd;
aud[1540]=16'h231;
aud[1541]=16'h28c;
aud[1542]=16'h2db;
aud[1543]=16'h31e;
aud[1544]=16'h353;
aud[1545]=16'h37a;
aud[1546]=16'h392;
aud[1547]=16'h39a;
aud[1548]=16'h392;
aud[1549]=16'h37a;
aud[1550]=16'h353;
aud[1551]=16'h31e;
aud[1552]=16'h2db;
aud[1553]=16'h28c;
aud[1554]=16'h231;
aud[1555]=16'h1cd;
aud[1556]=16'h161;
aud[1557]=16'hef;
aud[1558]=16'h78;
aud[1559]=16'h0;
aud[1560]=16'hff88;
aud[1561]=16'hff11;
aud[1562]=16'hfe9f;
aud[1563]=16'hfe33;
aud[1564]=16'hfdcf;
aud[1565]=16'hfd74;
aud[1566]=16'hfd25;
aud[1567]=16'hfce2;
aud[1568]=16'hfcad;
aud[1569]=16'hfc86;
aud[1570]=16'hfc6e;
aud[1571]=16'hfc66;
aud[1572]=16'hfc6e;
aud[1573]=16'hfc86;
aud[1574]=16'hfcad;
aud[1575]=16'hfce2;
aud[1576]=16'hfd25;
aud[1577]=16'hfd74;
aud[1578]=16'hfdcf;
aud[1579]=16'hfe33;
aud[1580]=16'hfe9f;
aud[1581]=16'hff11;
aud[1582]=16'hff88;
aud[1583]=16'h0;
aud[1584]=16'h78;
aud[1585]=16'hef;
aud[1586]=16'h161;
aud[1587]=16'h1cd;
aud[1588]=16'h231;
aud[1589]=16'h28c;
aud[1590]=16'h2db;
aud[1591]=16'h31e;
aud[1592]=16'h353;
aud[1593]=16'h37a;
aud[1594]=16'h392;
aud[1595]=16'h39a;
aud[1596]=16'h392;
aud[1597]=16'h37a;
aud[1598]=16'h353;
aud[1599]=16'h31e;
aud[1600]=16'h2db;
aud[1601]=16'h28c;
aud[1602]=16'h231;
aud[1603]=16'h1cd;
aud[1604]=16'h161;
aud[1605]=16'hef;
aud[1606]=16'h78;
aud[1607]=16'h0;
aud[1608]=16'hff88;
aud[1609]=16'hff11;
aud[1610]=16'hfe9f;
aud[1611]=16'hfe33;
aud[1612]=16'hfdcf;
aud[1613]=16'hfd74;
aud[1614]=16'hfd25;
aud[1615]=16'hfce2;
aud[1616]=16'hfcad;
aud[1617]=16'hfc86;
aud[1618]=16'hfc6e;
aud[1619]=16'hfc66;
aud[1620]=16'hfc6e;
aud[1621]=16'hfc86;
aud[1622]=16'hfcad;
aud[1623]=16'hfce2;
aud[1624]=16'hfd25;
aud[1625]=16'hfd74;
aud[1626]=16'hfdcf;
aud[1627]=16'hfe33;
aud[1628]=16'hfe9f;
aud[1629]=16'hff11;
aud[1630]=16'hff88;
aud[1631]=16'h0;
aud[1632]=16'h78;
aud[1633]=16'hef;
aud[1634]=16'h161;
aud[1635]=16'h1cd;
aud[1636]=16'h231;
aud[1637]=16'h28c;
aud[1638]=16'h2db;
aud[1639]=16'h31e;
aud[1640]=16'h353;
aud[1641]=16'h37a;
aud[1642]=16'h392;
aud[1643]=16'h39a;
aud[1644]=16'h392;
aud[1645]=16'h37a;
aud[1646]=16'h353;
aud[1647]=16'h31e;
aud[1648]=16'h2db;
aud[1649]=16'h28c;
aud[1650]=16'h231;
aud[1651]=16'h1cd;
aud[1652]=16'h161;
aud[1653]=16'hef;
aud[1654]=16'h78;
aud[1655]=16'h0;
aud[1656]=16'hff88;
aud[1657]=16'hff11;
aud[1658]=16'hfe9f;
aud[1659]=16'hfe33;
aud[1660]=16'hfdcf;
aud[1661]=16'hfd74;
aud[1662]=16'hfd25;
aud[1663]=16'hfce2;
aud[1664]=16'hfcad;
aud[1665]=16'hfc86;
aud[1666]=16'hfc6e;
aud[1667]=16'hfc66;
aud[1668]=16'hfc6e;
aud[1669]=16'hfc86;
aud[1670]=16'hfcad;
aud[1671]=16'hfce2;
aud[1672]=16'hfd25;
aud[1673]=16'hfd74;
aud[1674]=16'hfdcf;
aud[1675]=16'hfe33;
aud[1676]=16'hfe9f;
aud[1677]=16'hff11;
aud[1678]=16'hff88;
aud[1679]=16'h0;
aud[1680]=16'h78;
aud[1681]=16'hef;
aud[1682]=16'h161;
aud[1683]=16'h1cd;
aud[1684]=16'h231;
aud[1685]=16'h28c;
aud[1686]=16'h2db;
aud[1687]=16'h31e;
aud[1688]=16'h353;
aud[1689]=16'h37a;
aud[1690]=16'h392;
aud[1691]=16'h39a;
aud[1692]=16'h392;
aud[1693]=16'h37a;
aud[1694]=16'h353;
aud[1695]=16'h31e;
aud[1696]=16'h2db;
aud[1697]=16'h28c;
aud[1698]=16'h231;
aud[1699]=16'h1cd;
aud[1700]=16'h161;
aud[1701]=16'hef;
aud[1702]=16'h78;
aud[1703]=16'h0;
aud[1704]=16'hff88;
aud[1705]=16'hff11;
aud[1706]=16'hfe9f;
aud[1707]=16'hfe33;
aud[1708]=16'hfdcf;
aud[1709]=16'hfd74;
aud[1710]=16'hfd25;
aud[1711]=16'hfce2;
aud[1712]=16'hfcad;
aud[1713]=16'hfc86;
aud[1714]=16'hfc6e;
aud[1715]=16'hfc66;
aud[1716]=16'hfc6e;
aud[1717]=16'hfc86;
aud[1718]=16'hfcad;
aud[1719]=16'hfce2;
aud[1720]=16'hfd25;
aud[1721]=16'hfd74;
aud[1722]=16'hfdcf;
aud[1723]=16'hfe33;
aud[1724]=16'hfe9f;
aud[1725]=16'hff11;
aud[1726]=16'hff88;
aud[1727]=16'h0;
aud[1728]=16'h78;
aud[1729]=16'hef;
aud[1730]=16'h161;
aud[1731]=16'h1cd;
aud[1732]=16'h231;
aud[1733]=16'h28c;
aud[1734]=16'h2db;
aud[1735]=16'h31e;
aud[1736]=16'h353;
aud[1737]=16'h37a;
aud[1738]=16'h392;
aud[1739]=16'h39a;
aud[1740]=16'h392;
aud[1741]=16'h37a;
aud[1742]=16'h353;
aud[1743]=16'h31e;
aud[1744]=16'h2db;
aud[1745]=16'h28c;
aud[1746]=16'h231;
aud[1747]=16'h1cd;
aud[1748]=16'h161;
aud[1749]=16'hef;
aud[1750]=16'h78;
aud[1751]=16'h0;
aud[1752]=16'hff88;
aud[1753]=16'hff11;
aud[1754]=16'hfe9f;
aud[1755]=16'hfe33;
aud[1756]=16'hfdcf;
aud[1757]=16'hfd74;
aud[1758]=16'hfd25;
aud[1759]=16'hfce2;
aud[1760]=16'hfcad;
aud[1761]=16'hfc86;
aud[1762]=16'hfc6e;
aud[1763]=16'hfc66;
aud[1764]=16'hfc6e;
aud[1765]=16'hfc86;
aud[1766]=16'hfcad;
aud[1767]=16'hfce2;
aud[1768]=16'hfd25;
aud[1769]=16'hfd74;
aud[1770]=16'hfdcf;
aud[1771]=16'hfe33;
aud[1772]=16'hfe9f;
aud[1773]=16'hff11;
aud[1774]=16'hff88;
aud[1775]=16'h0;
aud[1776]=16'h78;
aud[1777]=16'hef;
aud[1778]=16'h161;
aud[1779]=16'h1cd;
aud[1780]=16'h231;
aud[1781]=16'h28c;
aud[1782]=16'h2db;
aud[1783]=16'h31e;
aud[1784]=16'h353;
aud[1785]=16'h37a;
aud[1786]=16'h392;
aud[1787]=16'h39a;
aud[1788]=16'h392;
aud[1789]=16'h37a;
aud[1790]=16'h353;
aud[1791]=16'h31e;
aud[1792]=16'h2db;
aud[1793]=16'h28c;
aud[1794]=16'h231;
aud[1795]=16'h1cd;
aud[1796]=16'h161;
aud[1797]=16'hef;
aud[1798]=16'h78;
aud[1799]=16'h0;
aud[1800]=16'hff88;
aud[1801]=16'hff11;
aud[1802]=16'hfe9f;
aud[1803]=16'hfe33;
aud[1804]=16'hfdcf;
aud[1805]=16'hfd74;
aud[1806]=16'hfd25;
aud[1807]=16'hfce2;
aud[1808]=16'hfcad;
aud[1809]=16'hfc86;
aud[1810]=16'hfc6e;
aud[1811]=16'hfc66;
aud[1812]=16'hfc6e;
aud[1813]=16'hfc86;
aud[1814]=16'hfcad;
aud[1815]=16'hfce2;
aud[1816]=16'hfd25;
aud[1817]=16'hfd74;
aud[1818]=16'hfdcf;
aud[1819]=16'hfe33;
aud[1820]=16'hfe9f;
aud[1821]=16'hff11;
aud[1822]=16'hff88;
aud[1823]=16'h0;
aud[1824]=16'h78;
aud[1825]=16'hef;
aud[1826]=16'h161;
aud[1827]=16'h1cd;
aud[1828]=16'h231;
aud[1829]=16'h28c;
aud[1830]=16'h2db;
aud[1831]=16'h31e;
aud[1832]=16'h353;
aud[1833]=16'h37a;
aud[1834]=16'h392;
aud[1835]=16'h39a;
aud[1836]=16'h392;
aud[1837]=16'h37a;
aud[1838]=16'h353;
aud[1839]=16'h31e;
aud[1840]=16'h2db;
aud[1841]=16'h28c;
aud[1842]=16'h231;
aud[1843]=16'h1cd;
aud[1844]=16'h161;
aud[1845]=16'hef;
aud[1846]=16'h78;
aud[1847]=16'h0;
aud[1848]=16'hff88;
aud[1849]=16'hff11;
aud[1850]=16'hfe9f;
aud[1851]=16'hfe33;
aud[1852]=16'hfdcf;
aud[1853]=16'hfd74;
aud[1854]=16'hfd25;
aud[1855]=16'hfce2;
aud[1856]=16'hfcad;
aud[1857]=16'hfc86;
aud[1858]=16'hfc6e;
aud[1859]=16'hfc66;
aud[1860]=16'hfc6e;
aud[1861]=16'hfc86;
aud[1862]=16'hfcad;
aud[1863]=16'hfce2;
aud[1864]=16'hfd25;
aud[1865]=16'hfd74;
aud[1866]=16'hfdcf;
aud[1867]=16'hfe33;
aud[1868]=16'hfe9f;
aud[1869]=16'hff11;
aud[1870]=16'hff88;
aud[1871]=16'h0;
aud[1872]=16'h78;
aud[1873]=16'hef;
aud[1874]=16'h161;
aud[1875]=16'h1cd;
aud[1876]=16'h231;
aud[1877]=16'h28c;
aud[1878]=16'h2db;
aud[1879]=16'h31e;
aud[1880]=16'h353;
aud[1881]=16'h37a;
aud[1882]=16'h392;
aud[1883]=16'h39a;
aud[1884]=16'h392;
aud[1885]=16'h37a;
aud[1886]=16'h353;
aud[1887]=16'h31e;
aud[1888]=16'h2db;
aud[1889]=16'h28c;
aud[1890]=16'h231;
aud[1891]=16'h1cd;
aud[1892]=16'h161;
aud[1893]=16'hef;
aud[1894]=16'h78;
aud[1895]=16'h0;
aud[1896]=16'hff88;
aud[1897]=16'hff11;
aud[1898]=16'hfe9f;
aud[1899]=16'hfe33;
aud[1900]=16'hfdcf;
aud[1901]=16'hfd74;
aud[1902]=16'hfd25;
aud[1903]=16'hfce2;
aud[1904]=16'hfcad;
aud[1905]=16'hfc86;
aud[1906]=16'hfc6e;
aud[1907]=16'hfc66;
aud[1908]=16'hfc6e;
aud[1909]=16'hfc86;
aud[1910]=16'hfcad;
aud[1911]=16'hfce2;
aud[1912]=16'hfd25;
aud[1913]=16'hfd74;
aud[1914]=16'hfdcf;
aud[1915]=16'hfe33;
aud[1916]=16'hfe9f;
aud[1917]=16'hff11;
aud[1918]=16'hff88;
aud[1919]=16'h0;
aud[1920]=16'h78;
aud[1921]=16'hef;
aud[1922]=16'h161;
aud[1923]=16'h1cd;
aud[1924]=16'h231;
aud[1925]=16'h28c;
aud[1926]=16'h2db;
aud[1927]=16'h31e;
aud[1928]=16'h353;
aud[1929]=16'h37a;
aud[1930]=16'h392;
aud[1931]=16'h39a;
aud[1932]=16'h392;
aud[1933]=16'h37a;
aud[1934]=16'h353;
aud[1935]=16'h31e;
aud[1936]=16'h2db;
aud[1937]=16'h28c;
aud[1938]=16'h231;
aud[1939]=16'h1cd;
aud[1940]=16'h161;
aud[1941]=16'hef;
aud[1942]=16'h78;
aud[1943]=16'h0;
aud[1944]=16'hff88;
aud[1945]=16'hff11;
aud[1946]=16'hfe9f;
aud[1947]=16'hfe33;
aud[1948]=16'hfdcf;
aud[1949]=16'hfd74;
aud[1950]=16'hfd25;
aud[1951]=16'hfce2;
aud[1952]=16'hfcad;
aud[1953]=16'hfc86;
aud[1954]=16'hfc6e;
aud[1955]=16'hfc66;
aud[1956]=16'hfc6e;
aud[1957]=16'hfc86;
aud[1958]=16'hfcad;
aud[1959]=16'hfce2;
aud[1960]=16'hfd25;
aud[1961]=16'hfd74;
aud[1962]=16'hfdcf;
aud[1963]=16'hfe33;
aud[1964]=16'hfe9f;
aud[1965]=16'hff11;
aud[1966]=16'hff88;
aud[1967]=16'h0;
aud[1968]=16'h78;
aud[1969]=16'hef;
aud[1970]=16'h161;
aud[1971]=16'h1cd;
aud[1972]=16'h231;
aud[1973]=16'h28c;
aud[1974]=16'h2db;
aud[1975]=16'h31e;
aud[1976]=16'h353;
aud[1977]=16'h37a;
aud[1978]=16'h392;
aud[1979]=16'h39a;
aud[1980]=16'h392;
aud[1981]=16'h37a;
aud[1982]=16'h353;
aud[1983]=16'h31e;
aud[1984]=16'h2db;
aud[1985]=16'h28c;
aud[1986]=16'h231;
aud[1987]=16'h1cd;
aud[1988]=16'h161;
aud[1989]=16'hef;
aud[1990]=16'h78;
aud[1991]=16'h0;
aud[1992]=16'hff88;
aud[1993]=16'hff11;
aud[1994]=16'hfe9f;
aud[1995]=16'hfe33;
aud[1996]=16'hfdcf;
aud[1997]=16'hfd74;
aud[1998]=16'hfd25;
aud[1999]=16'hfce2;

end


endmodule